library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cv17_36 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cv17_36 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"C3",X"D9",X"0A",X"00",X"00",X"F5",X"C5",X"D5",X"E5",X"C3",X"88",X"00",X"00",
		X"F5",X"C5",X"D5",X"E5",X"3E",X"80",X"32",X"72",X"20",X"21",X"C0",X"20",X"35",X"CD",X"DD",X"17",
		X"DB",X"01",X"0F",X"DA",X"67",X"00",X"3A",X"EA",X"20",X"A7",X"CA",X"42",X"00",X"3A",X"EB",X"20",
		X"FE",X"99",X"CA",X"3E",X"00",X"C6",X"01",X"27",X"32",X"EB",X"20",X"CD",X"2E",X"19",X"AF",X"32",
		X"EA",X"20",X"3A",X"E9",X"20",X"A7",X"CA",X"82",X"00",X"3A",X"EF",X"20",X"A7",X"C2",X"6F",X"00",
		X"3A",X"EB",X"20",X"A7",X"C2",X"5D",X"00",X"CD",X"AE",X"0A",X"C3",X"82",X"00",X"3A",X"93",X"20",
		X"A7",X"C2",X"82",X"00",X"C3",X"4C",X"07",X"3E",X"01",X"32",X"EA",X"20",X"C3",X"3F",X"00",X"CD",
		X"5C",X"17",X"3A",X"32",X"20",X"32",X"80",X"20",X"CD",X"E3",X"00",X"CD",X"30",X"02",X"CD",X"FF",
		X"08",X"00",X"E1",X"D1",X"C1",X"F1",X"FB",X"C9",X"AF",X"32",X"72",X"20",X"3A",X"E9",X"20",X"A7",
		X"CA",X"82",X"00",X"3A",X"EF",X"20",X"A7",X"C2",X"A1",X"00",X"3A",X"C1",X"20",X"0F",X"D2",X"82",
		X"00",X"21",X"20",X"20",X"CD",X"33",X"02",X"CD",X"24",X"01",X"C3",X"82",X"00",X"CD",X"6A",X"08",
		X"E5",X"7E",X"23",X"66",X"6F",X"22",X"09",X"20",X"22",X"0B",X"20",X"E1",X"2B",X"7E",X"FE",X"03",
		X"C2",X"C4",X"00",X"3D",X"32",X"08",X"20",X"FE",X"FE",X"3E",X"00",X"C2",X"CF",X"00",X"3C",X"32",
		X"0D",X"20",X"C9",X"EB",X"6E",X"26",X"00",X"79",X"B7",X"CA",X"E1",X"00",X"29",X"3D",X"C2",X"DC",
		X"00",X"EB",X"C9",X"21",X"02",X"20",X"7E",X"A7",X"C2",X"09",X"15",X"E5",X"3A",X"06",X"20",X"6F",
		X"3A",X"67",X"20",X"67",X"7E",X"A7",X"E1",X"CA",X"19",X"01",X"23",X"23",X"7E",X"23",X"46",X"E6",
		X"FE",X"07",X"07",X"07",X"5F",X"16",X"00",X"21",X"00",X"1C",X"19",X"EB",X"78",X"A7",X"C4",X"1E",
		X"01",X"2A",X"0B",X"20",X"06",X"10",X"CD",X"F5",X"15",X"AF",X"32",X"00",X"20",X"C9",X"21",X"30",
		X"00",X"19",X"EB",X"C9",X"3A",X"68",X"20",X"A7",X"C8",X"3A",X"00",X"20",X"A7",X"C0",X"3A",X"67",
		X"20",X"67",X"3A",X"06",X"20",X"16",X"02",X"3C",X"FE",X"37",X"CC",X"84",X"01",X"6F",X"46",X"05",
		X"C2",X"37",X"01",X"32",X"06",X"20",X"CD",X"5D",X"01",X"61",X"22",X"0B",X"20",X"7D",X"FE",X"28",
		X"DA",X"58",X"19",X"7A",X"32",X"04",X"20",X"3E",X"01",X"32",X"00",X"20",X"C9",X"16",X"00",X"7D",
		X"21",X"09",X"20",X"46",X"23",X"4E",X"FE",X"0B",X"FA",X"77",X"01",X"DE",X"0B",X"5F",X"78",X"C6",
		X"10",X"47",X"7B",X"14",X"C3",X"66",X"01",X"68",X"A7",X"C8",X"5F",X"79",X"C6",X"10",X"4F",X"7B",
		X"3D",X"C3",X"78",X"01",X"15",X"CA",X"B5",X"01",X"21",X"06",X"20",X"36",X"00",X"23",X"4E",X"36",
		X"00",X"CD",X"C1",X"01",X"21",X"05",X"20",X"7E",X"3C",X"E6",X"01",X"77",X"AF",X"21",X"67",X"20",
		X"66",X"C9",X"21",X"00",X"22",X"C3",X"AB",X"01",X"21",X"00",X"21",X"06",X"37",X"36",X"01",X"23",
		X"05",X"C2",X"AD",X"01",X"C9",X"E1",X"C9",X"3E",X"01",X"06",X"E0",X"21",X"02",X"24",X"C3",X"85",
		X"14",X"23",X"46",X"23",X"79",X"86",X"77",X"23",X"78",X"86",X"77",X"C9",X"06",X"C0",X"11",X"00",
		X"1B",X"21",X"00",X"20",X"C3",X"14",X"1A",X"21",X"42",X"21",X"C3",X"E0",X"01",X"21",X"42",X"22",
		X"0E",X"04",X"11",X"20",X"1D",X"D5",X"06",X"2C",X"CD",X"14",X"1A",X"D1",X"0D",X"C2",X"E5",X"01",
		X"C9",X"3E",X"01",X"C3",X"03",X"02",X"3E",X"01",X"C3",X"FC",X"01",X"AF",X"11",X"42",X"22",X"C3",
		X"06",X"02",X"AF",X"11",X"42",X"21",X"32",X"81",X"20",X"01",X"02",X"16",X"21",X"06",X"28",X"3E",
		X"04",X"F5",X"C5",X"3A",X"81",X"20",X"A7",X"C2",X"2A",X"02",X"CD",X"4F",X"1A",X"C1",X"F1",X"3D",
		X"C8",X"D5",X"11",X"E0",X"02",X"19",X"D1",X"C3",X"11",X"02",X"CD",X"46",X"14",X"C3",X"1D",X"02",
		X"21",X"10",X"20",X"7E",X"FE",X"FF",X"C8",X"FE",X"FE",X"CA",X"69",X"02",X"23",X"46",X"4F",X"B0",
		X"79",X"C2",X"5F",X"02",X"23",X"7E",X"A7",X"C2",X"70",X"02",X"23",X"5E",X"23",X"56",X"E5",X"EB",
		X"E5",X"21",X"57",X"02",X"E3",X"D5",X"E9",X"E1",X"11",X"0C",X"00",X"19",X"C3",X"33",X"02",X"05",
		X"04",X"C2",X"65",X"02",X"3D",X"05",X"70",X"2B",X"77",X"11",X"10",X"00",X"19",X"C3",X"33",X"02",
		X"35",X"2B",X"2B",X"C3",X"69",X"02",X"E1",X"23",X"7E",X"FE",X"FF",X"CA",X"2C",X"03",X"23",X"35",
		X"C0",X"47",X"AF",X"32",X"68",X"20",X"32",X"69",X"20",X"3E",X"30",X"32",X"6A",X"20",X"78",X"36",
		X"05",X"23",X"35",X"C2",X"8B",X"03",X"2A",X"1A",X"20",X"06",X"10",X"CD",X"00",X"14",X"21",X"10",
		X"20",X"11",X"10",X"1B",X"06",X"10",X"CD",X"14",X"1A",X"06",X"00",X"CD",X"BE",X"19",X"3A",X"6D",
		X"20",X"A7",X"C0",X"3A",X"EF",X"20",X"A7",X"C8",X"31",X"00",X"24",X"FB",X"CD",X"BA",X"19",X"CD",
		X"1A",X"09",X"A7",X"CA",X"80",X"16",X"CD",X"DD",X"18",X"7E",X"A7",X"CA",X"20",X"03",X"3A",X"CE",
		X"20",X"A7",X"CA",X"20",X"03",X"3A",X"67",X"20",X"F5",X"0F",X"DA",X"26",X"03",X"CD",X"F6",X"01",
		X"CD",X"5F",X"08",X"73",X"23",X"72",X"2B",X"2B",X"70",X"CD",X"CC",X"01",X"F1",X"0F",X"3E",X"21",
		X"06",X"00",X"D2",X"F9",X"02",X"06",X"20",X"3E",X"22",X"32",X"67",X"20",X"CD",X"A5",X"0A",X"AF",
		X"32",X"11",X"20",X"F3",X"78",X"D3",X"05",X"01",X"0A",X"00",X"05",X"C2",X"0A",X"03",X"0D",X"C2",
		X"0A",X"03",X"FB",X"3C",X"32",X"98",X"20",X"CD",X"C5",X"09",X"CD",X"65",X"1A",X"C3",X"E3",X"07",
		X"CD",X"65",X"1A",X"C3",X"01",X"08",X"CD",X"F1",X"01",X"C3",X"E0",X"02",X"21",X"68",X"20",X"36",
		X"01",X"23",X"7E",X"A7",X"C3",X"A0",X"03",X"2B",X"36",X"01",X"3A",X"1B",X"20",X"47",X"3A",X"EF",
		X"20",X"A7",X"C2",X"53",X"03",X"3A",X"1D",X"20",X"0F",X"DA",X"71",X"03",X"0F",X"DA",X"7E",X"03",
		X"C3",X"5F",X"03",X"CD",X"D0",X"17",X"07",X"07",X"DA",X"71",X"03",X"07",X"DA",X"7E",X"03",X"21",
		X"18",X"20",X"CD",X"1D",X"1A",X"CD",X"2D",X"1A",X"CD",X"15",X"14",X"3E",X"00",X"32",X"12",X"20",
		X"C9",X"78",X"FE",X"D9",X"CA",X"5F",X"03",X"3C",X"32",X"1B",X"20",X"C3",X"5F",X"03",X"78",X"FE",
		X"30",X"CA",X"5F",X"03",X"3D",X"32",X"1B",X"20",X"C3",X"5F",X"03",X"3C",X"E6",X"01",X"32",X"15",
		X"20",X"07",X"07",X"07",X"07",X"21",X"70",X"1C",X"85",X"6F",X"22",X"18",X"20",X"C3",X"5F",X"03",
		X"C2",X"3A",X"03",X"23",X"35",X"C2",X"3A",X"03",X"C3",X"37",X"03",X"11",X"2A",X"20",X"CD",X"E8",
		X"19",X"E1",X"D0",X"23",X"7E",X"A7",X"C8",X"FE",X"01",X"CA",X"EA",X"03",X"FE",X"02",X"CA",X"FA",
		X"03",X"23",X"FE",X"03",X"C2",X"1A",X"04",X"35",X"CA",X"26",X"04",X"7E",X"FE",X"0F",X"C0",X"E5",
		X"CD",X"20",X"04",X"CD",X"24",X"15",X"E1",X"23",X"34",X"23",X"23",X"35",X"35",X"23",X"35",X"35",
		X"35",X"23",X"36",X"08",X"CD",X"20",X"04",X"C3",X"23",X"14",X"3C",X"77",X"3A",X"1B",X"20",X"C6",
		X"08",X"32",X"2A",X"20",X"CD",X"20",X"04",X"C3",X"23",X"14",X"CD",X"20",X"04",X"D5",X"E5",X"C5",
		X"CD",X"24",X"15",X"C1",X"E1",X"D1",X"3A",X"2C",X"20",X"85",X"6F",X"32",X"29",X"20",X"CD",X"C0",
		X"15",X"3A",X"61",X"20",X"A7",X"C8",X"32",X"02",X"20",X"C9",X"FE",X"05",X"C8",X"C3",X"26",X"04",
		X"21",X"27",X"20",X"C3",X"1D",X"1A",X"CD",X"20",X"04",X"CD",X"24",X"15",X"21",X"25",X"20",X"11",
		X"25",X"1B",X"06",X"07",X"CD",X"14",X"1A",X"2A",X"8D",X"20",X"2C",X"7D",X"FE",X"63",X"DA",X"43",
		X"04",X"2E",X"54",X"22",X"8D",X"20",X"2A",X"8F",X"20",X"2C",X"22",X"8F",X"20",X"3A",X"84",X"20",
		X"A7",X"C0",X"7E",X"E6",X"01",X"01",X"29",X"02",X"C2",X"5E",X"04",X"01",X"E0",X"FE",X"21",X"8A",
		X"20",X"71",X"23",X"23",X"70",X"C9",X"E1",X"3A",X"32",X"1B",X"32",X"32",X"20",X"2A",X"38",X"20",
		X"7D",X"B4",X"C2",X"7A",X"04",X"2B",X"22",X"38",X"20",X"C9",X"11",X"35",X"20",X"3E",X"F9",X"CD",
		X"40",X"05",X"3A",X"46",X"20",X"32",X"70",X"20",X"3A",X"56",X"20",X"32",X"71",X"20",X"CD",X"53",
		X"05",X"3A",X"78",X"20",X"A7",X"21",X"35",X"20",X"C2",X"4B",X"05",X"11",X"30",X"1B",X"21",X"30",
		X"20",X"06",X"10",X"C3",X"14",X"1A",X"E1",X"3A",X"6E",X"20",X"A7",X"C0",X"3A",X"80",X"20",X"FE",
		X"01",X"C0",X"11",X"45",X"20",X"3E",X"ED",X"CD",X"40",X"05",X"3A",X"36",X"20",X"32",X"70",X"20",
		X"3A",X"56",X"20",X"32",X"71",X"20",X"CD",X"53",X"05",X"3A",X"76",X"20",X"FE",X"10",X"DA",X"D7",
		X"04",X"3A",X"48",X"1B",X"32",X"76",X"20",X"3A",X"78",X"20",X"A7",X"21",X"45",X"20",X"C2",X"4B",
		X"05",X"11",X"40",X"1B",X"21",X"40",X"20",X"06",X"10",X"CD",X"14",X"1A",X"3A",X"82",X"20",X"3D",
		X"C2",X"F8",X"04",X"3E",X"01",X"32",X"6E",X"20",X"2A",X"76",X"20",X"C3",X"6C",X"06",X"E1",X"11",
		X"55",X"20",X"3E",X"DB",X"CD",X"40",X"05",X"3A",X"46",X"20",X"32",X"70",X"20",X"3A",X"36",X"20",
		X"32",X"71",X"20",X"CD",X"53",X"05",X"3A",X"76",X"20",X"FE",X"15",X"DA",X"24",X"05",X"3A",X"58",
		X"1B",X"32",X"76",X"20",X"3A",X"78",X"20",X"A7",X"21",X"55",X"20",X"C2",X"4B",X"05",X"11",X"50",
		X"1B",X"21",X"50",X"20",X"06",X"10",X"CD",X"14",X"1A",X"2A",X"76",X"20",X"22",X"58",X"20",X"C9",
		X"32",X"7F",X"20",X"21",X"73",X"20",X"06",X"0B",X"C3",X"14",X"1A",X"11",X"73",X"20",X"06",X"0B",
		X"C3",X"14",X"1A",X"21",X"73",X"20",X"7E",X"E6",X"80",X"C2",X"B0",X"05",X"3A",X"C1",X"20",X"FE",
		X"04",X"3A",X"69",X"20",X"CA",X"A6",X"05",X"A7",X"C8",X"23",X"36",X"00",X"3A",X"70",X"20",X"A7",
		X"CA",X"79",X"05",X"47",X"3A",X"CF",X"20",X"B8",X"D0",X"3A",X"71",X"20",X"A7",X"CA",X"86",X"05",
		X"47",X"3A",X"CF",X"20",X"B8",X"D0",X"23",X"7E",X"A7",X"CA",X"09",X"06",X"2A",X"76",X"20",X"4E",
		X"23",X"22",X"76",X"20",X"CD",X"1D",X"06",X"D0",X"CD",X"5D",X"01",X"79",X"C6",X"07",X"67",X"7D",
		X"D6",X"0A",X"6F",X"22",X"7B",X"20",X"21",X"73",X"20",X"7E",X"F6",X"80",X"77",X"23",X"34",X"C9",
		X"11",X"7C",X"20",X"CD",X"E8",X"19",X"D0",X"23",X"7E",X"E6",X"01",X"C2",X"32",X"06",X"23",X"34",
		X"CD",X"63",X"06",X"3A",X"79",X"20",X"C6",X"03",X"21",X"7F",X"20",X"BE",X"DA",X"D1",X"05",X"D6",
		X"0C",X"32",X"79",X"20",X"3A",X"7B",X"20",X"47",X"3A",X"7E",X"20",X"80",X"32",X"7B",X"20",X"CD",
		X"5A",X"06",X"3A",X"7B",X"20",X"FE",X"15",X"DA",X"00",X"06",X"3A",X"61",X"20",X"A7",X"C8",X"3A",
		X"7B",X"20",X"FE",X"1E",X"DA",X"00",X"06",X"FE",X"27",X"D2",X"00",X"06",X"97",X"32",X"15",X"20",
		X"3A",X"73",X"20",X"F6",X"01",X"32",X"73",X"20",X"C9",X"3A",X"1B",X"20",X"C6",X"08",X"67",X"CD",
		X"5A",X"15",X"79",X"FE",X"0C",X"DA",X"94",X"05",X"0E",X"0B",X"C3",X"94",X"05",X"0D",X"3A",X"67",
		X"20",X"67",X"69",X"16",X"05",X"7E",X"A7",X"37",X"C0",X"7D",X"C6",X"0B",X"6F",X"15",X"C2",X"25",
		X"06",X"C9",X"21",X"78",X"20",X"35",X"7E",X"FE",X"03",X"C2",X"55",X"06",X"CD",X"63",X"06",X"21",
		X"DC",X"1C",X"22",X"79",X"20",X"21",X"7C",X"20",X"35",X"35",X"2B",X"35",X"35",X"3E",X"06",X"32",
		X"7D",X"20",X"C3",X"5A",X"06",X"A7",X"C0",X"C3",X"63",X"06",X"21",X"79",X"20",X"CD",X"1D",X"1A",
		X"C3",X"C0",X"15",X"21",X"79",X"20",X"CD",X"1D",X"1A",X"C3",X"24",X"15",X"22",X"48",X"20",X"C9",
		X"E1",X"3A",X"80",X"20",X"FE",X"02",X"C0",X"21",X"83",X"20",X"7E",X"A7",X"CA",X"FF",X"04",X"3A",
		X"56",X"20",X"A7",X"C2",X"FF",X"04",X"23",X"7E",X"A7",X"C2",X"99",X"06",X"3A",X"82",X"20",X"FE",
		X"08",X"DA",X"FF",X"04",X"36",X"01",X"CD",X"23",X"07",X"11",X"8A",X"20",X"CD",X"E8",X"19",X"D0",
		X"21",X"85",X"20",X"7E",X"A7",X"C2",X"C4",X"06",X"21",X"8A",X"20",X"7E",X"23",X"23",X"86",X"32",
		X"8A",X"20",X"CD",X"23",X"07",X"21",X"8A",X"20",X"7E",X"FE",X"28",X"DA",X"E4",X"06",X"FE",X"E1",
		X"D2",X"E4",X"06",X"C9",X"06",X"FE",X"CD",X"BE",X"19",X"23",X"35",X"7E",X"FE",X"1F",X"CA",X"32",
		X"07",X"FE",X"18",X"CA",X"F7",X"06",X"A7",X"C0",X"06",X"EF",X"21",X"98",X"20",X"7E",X"A0",X"77",
		X"E6",X"20",X"D3",X"05",X"CD",X"29",X"07",X"CD",X"84",X"14",X"21",X"83",X"20",X"06",X"0A",X"CD",
		X"46",X"07",X"06",X"FE",X"C3",X"BE",X"19",X"3E",X"01",X"32",X"F1",X"20",X"2A",X"8D",X"20",X"46",
		X"0E",X"04",X"21",X"50",X"1D",X"11",X"4C",X"1D",X"1A",X"B8",X"CA",X"13",X"07",X"23",X"13",X"0D",
		X"C2",X"08",X"07",X"7E",X"32",X"87",X"20",X"26",X"00",X"68",X"22",X"F2",X"20",X"CD",X"29",X"07",
		X"C3",X"DD",X"08",X"CD",X"29",X"07",X"C3",X"15",X"14",X"21",X"87",X"20",X"CD",X"1D",X"1A",X"C3",
		X"2D",X"1A",X"06",X"10",X"21",X"98",X"20",X"7E",X"B0",X"77",X"CD",X"8C",X"17",X"21",X"7C",X"1D",
		X"22",X"87",X"20",X"C3",X"23",X"07",X"11",X"83",X"1B",X"C3",X"14",X"1A",X"3E",X"01",X"32",X"93",
		X"20",X"31",X"00",X"24",X"FB",X"CD",X"60",X"19",X"CD",X"C5",X"09",X"21",X"13",X"30",X"11",X"F3",
		X"1F",X"0E",X"04",X"CD",X"DF",X"08",X"3A",X"EB",X"20",X"3D",X"21",X"10",X"28",X"0E",X"14",X"C2",
		X"3E",X"08",X"11",X"CF",X"1A",X"CD",X"DF",X"08",X"DB",X"01",X"E6",X"04",X"CA",X"66",X"07",X"06",
		X"99",X"AF",X"32",X"CE",X"20",X"3A",X"EB",X"20",X"80",X"27",X"32",X"EB",X"20",X"CD",X"2E",X"19",
		X"21",X"00",X"00",X"22",X"F8",X"20",X"22",X"FC",X"20",X"CD",X"0F",X"19",X"CD",X"15",X"19",X"CD",
		X"BA",X"19",X"21",X"01",X"01",X"7C",X"32",X"EF",X"20",X"22",X"E7",X"20",X"22",X"E5",X"20",X"CD",
		X"3D",X"19",X"CD",X"D7",X"01",X"CD",X"DD",X"01",X"CD",X"B5",X"08",X"32",X"FF",X"21",X"32",X"FF",
		X"22",X"CD",X"C8",X"08",X"AF",X"32",X"FE",X"21",X"32",X"FE",X"22",X"CD",X"A8",X"01",X"CD",X"A2",
		X"01",X"CD",X"5B",X"14",X"21",X"78",X"38",X"22",X"FC",X"21",X"22",X"FC",X"22",X"CD",X"CC",X"01",
		X"CD",X"65",X"1A",X"CD",X"71",X"08",X"CD",X"C5",X"09",X"00",X"AF",X"32",X"C1",X"20",X"CD",X"B7",
		X"01",X"3A",X"67",X"20",X"0F",X"DA",X"59",X"08",X"CD",X"FB",X"01",X"CD",X"B7",X"01",X"CD",X"AD");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
