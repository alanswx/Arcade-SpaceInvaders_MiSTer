library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cv19_34 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cv19_34 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CD",X"29",X"1A",X"C5",X"E5",X"AF",X"77",X"23",X"77",X"23",X"E1",X"01",X"20",X"00",X"09",X"C1",
		X"05",X"C2",X"03",X"14",X"C9",X"C5",X"1A",X"77",X"13",X"01",X"20",X"00",X"09",X"C1",X"05",X"C2",
		X"15",X"14",X"C9",X"CD",X"29",X"1A",X"D5",X"CD",X"D3",X"00",X"7B",X"B6",X"77",X"23",X"7A",X"B6",
		X"77",X"11",X"1F",X"00",X"19",X"D1",X"13",X"05",X"C2",X"26",X"14",X"C9",X"21",X"F3",X"76",X"22",
		X"00",X"20",X"21",X"00",X"20",X"E9",X"C5",X"E5",X"7E",X"12",X"13",X"23",X"0D",X"C2",X"48",X"14",
		X"E1",X"01",X"20",X"00",X"09",X"C1",X"05",X"C2",X"46",X"14",X"C9",X"21",X"00",X"00",X"06",X"02",
		X"11",X"A7",X"14",X"0E",X"0C",X"AF",X"86",X"CE",X"00",X"2C",X"C2",X"66",X"14",X"EB",X"BE",X"C4",
		X"3C",X"14",X"2B",X"EB",X"24",X"0D",X"C2",X"65",X"14",X"05",X"C8",X"0E",X"0B",X"3E",X"09",X"84",
		X"67",X"C3",X"65",X"14",X"AF",X"C5",X"77",X"01",X"20",X"00",X"09",X"C1",X"05",X"C2",X"85",X"14",
		X"C9",X"0E",X"13",X"2F",X"D9",X"30",X"A8",X"C1",X"2D",X"39",X"38",X"60",X"F4",X"A2",X"FC",X"9C",
		X"0D",X"C2",X"BF",X"0B",X"C6",X"7F",X"3D",X"1D",X"00",X"3A",X"25",X"20",X"FE",X"05",X"C8",X"FE",
		X"02",X"C0",X"3A",X"29",X"20",X"FE",X"D8",X"47",X"D2",X"01",X"15",X"3A",X"02",X"20",X"A7",X"C8",
		X"78",X"FE",X"CE",X"D2",X"64",X"15",X"C6",X"06",X"47",X"3A",X"09",X"20",X"FE",X"90",X"D2",X"D5",
		X"14",X"B8",X"D2",X"01",X"15",X"68",X"CD",X"4D",X"15",X"3A",X"2A",X"20",X"67",X"CD",X"5A",X"15",
		X"22",X"64",X"20",X"3E",X"05",X"32",X"25",X"20",X"CD",X"6C",X"15",X"7E",X"A7",X"CA",X"01",X"15",
		X"36",X"00",X"CD",X"4E",X"0A",X"CD",X"1D",X"1A",X"CD",X"F5",X"15",X"3E",X"10",X"32",X"03",X"20",
		X"C9",X"3E",X"03",X"32",X"25",X"20",X"C3",X"1B",X"15",X"21",X"03",X"20",X"35",X"C0",X"2A",X"64",
		X"20",X"06",X"10",X"CD",X"00",X"14",X"3E",X"04",X"32",X"25",X"20",X"AF",X"32",X"02",X"20",X"06",
		X"F7",X"C3",X"BE",X"19",X"CD",X"29",X"1A",X"D5",X"CD",X"D3",X"00",X"7B",X"2F",X"A6",X"77",X"23",
		X"7A",X"2F",X"A6",X"77",X"11",X"1F",X"00",X"19",X"D1",X"13",X"05",X"C2",X"27",X"15",X"C9",X"0E",
		X"00",X"BC",X"D4",X"7B",X"15",X"BC",X"D0",X"C6",X"10",X"0C",X"C3",X"45",X"15",X"3A",X"09",X"20",
		X"65",X"CD",X"3F",X"15",X"41",X"05",X"DE",X"10",X"6F",X"C9",X"3A",X"0A",X"20",X"CD",X"3F",X"15",
		X"DE",X"10",X"67",X"C9",X"3E",X"01",X"32",X"85",X"20",X"C3",X"16",X"15",X"78",X"07",X"07",X"07",
		X"80",X"80",X"80",X"81",X"3D",X"6F",X"3A",X"67",X"20",X"67",X"C9",X"0C",X"C6",X"10",X"FA",X"7B",
		X"15",X"C9",X"CD",X"A9",X"14",X"3A",X"0D",X"20",X"A7",X"C2",X"A5",X"15",X"21",X"A4",X"3E",X"CD",
		X"B3",X"15",X"D0",X"06",X"FE",X"3E",X"01",X"32",X"0D",X"20",X"78",X"32",X"08",X"20",X"3A",X"0E",
		X"20",X"32",X"07",X"20",X"C9",X"21",X"24",X"25",X"CD",X"B3",X"15",X"D0",X"CD",X"E7",X"18",X"AF",
		X"C3",X"97",X"15",X"06",X"17",X"7E",X"A7",X"37",X"C0",X"23",X"05",X"C2",X"B5",X"15",X"B7",X"C9",
		X"CD",X"29",X"1A",X"79",X"F5",X"0E",X"00",X"F1",X"F5",X"D5",X"C5",X"4F",X"CD",X"D3",X"00",X"C1",
		X"7B",X"A6",X"CA",X"D7",X"15",X"0E",X"01",X"7B",X"B6",X"77",X"23",X"7A",X"A6",X"CA",X"E2",X"15",
		X"0E",X"01",X"7A",X"B6",X"77",X"11",X"1F",X"00",X"19",X"D1",X"13",X"05",X"C2",X"C7",X"15",X"F1",
		X"79",X"32",X"61",X"20",X"C9",X"CD",X"2D",X"1A",X"C5",X"01",X"1F",X"00",X"1A",X"77",X"23",X"13",
		X"70",X"09",X"C1",X"05",X"C2",X"F8",X"15",X"C9",X"CD",X"26",X"16",X"01",X"00",X"37",X"7E",X"A7",
		X"CA",X"14",X"16",X"0C",X"23",X"05",X"C2",X"0E",X"16",X"79",X"32",X"82",X"20",X"FE",X"01",X"C0",
		X"21",X"6B",X"20",X"36",X"01",X"C9",X"2E",X"00",X"3A",X"67",X"20",X"67",X"C9",X"3A",X"15",X"20",
		X"FE",X"FF",X"C0",X"21",X"10",X"20",X"7E",X"23",X"46",X"B0",X"C0",X"3A",X"25",X"20",X"A7",X"C0",
		X"3A",X"EF",X"20",X"A7",X"CA",X"67",X"16",X"3A",X"2D",X"20",X"A7",X"C2",X"5D",X"16",X"CD",X"D0",
		X"17",X"E6",X"10",X"C8",X"3E",X"01",X"32",X"25",X"20",X"32",X"2D",X"20",X"C9",X"CD",X"D0",X"17",
		X"E6",X"10",X"C0",X"32",X"2D",X"20",X"C9",X"21",X"25",X"20",X"36",X"01",X"2A",X"ED",X"20",X"23",
		X"7D",X"FE",X"7E",X"DA",X"78",X"16",X"2E",X"74",X"22",X"ED",X"20",X"7E",X"32",X"1D",X"20",X"C9",
		X"AF",X"CD",X"71",X"1A",X"CD",X"FA",X"18",X"36",X"00",X"CD",X"B9",X"09",X"23",X"11",X"F5",X"20",
		X"1A",X"BE",X"1B",X"2B",X"1A",X"CA",X"9E",X"16",X"D2",X"AB",X"16",X"C3",X"A2",X"16",X"BE",X"D2",
		X"AB",X"16",X"7E",X"12",X"13",X"23",X"7E",X"12",X"CD",X"37",X"19",X"3A",X"CE",X"20",X"A7",X"CA",
		X"DC",X"16",X"21",X"03",X"28",X"11",X"A6",X"1A",X"0E",X"14",X"CD",X"82",X"0A",X"25",X"25",X"06",
		X"1B",X"3A",X"67",X"20",X"0F",X"DA",X"CA",X"16",X"06",X"1C",X"78",X"CD",X"EB",X"08",X"CD",X"A0",
		X"0A",X"CD",X"DD",X"18",X"7E",X"A7",X"CA",X"DC",X"16",X"C3",X"D5",X"02",X"21",X"18",X"2D",X"11",
		X"A6",X"1A",X"0E",X"0A",X"CD",X"82",X"0A",X"CD",X"A5",X"0A",X"CD",X"C5",X"09",X"AF",X"32",X"EF",
		X"20",X"D3",X"05",X"CD",X"B4",X"19",X"C3",X"88",X"0B",X"31",X"00",X"24",X"FB",X"AF",X"32",X"15",
		X"20",X"CD",X"A9",X"14",X"06",X"04",X"CD",X"F0",X"18",X"CD",X"48",X"0A",X"C2",X"01",X"17",X"CD",
		X"BA",X"19",X"21",X"01",X"27",X"CD",X"DC",X"19",X"AF",X"CD",X"71",X"1A",X"06",X"FB",X"C3",X"52",
		X"19",X"CD",X"3D",X"17",X"11",X"B8",X"1C",X"21",X"A1",X"1A",X"0E",X"04",X"47",X"1A",X"B8",X"D2",
		X"38",X"17",X"23",X"13",X"0D",X"C2",X"2D",X"17",X"7E",X"32",X"CF",X"20",X"C9",X"CD",X"B9",X"09",
		X"7E",X"23",X"66",X"6F",X"29",X"29",X"29",X"29",X"7C",X"C9",X"3A",X"25",X"20",X"FE",X"00",X"C2",
		X"57",X"17",X"06",X"FD",X"C3",X"BE",X"19",X"06",X"02",X"C3",X"F0",X"18",X"21",X"9B",X"20",X"35",
		X"CC",X"89",X"17",X"3A",X"68",X"20",X"A7",X"CA",X"89",X"17",X"21",X"96",X"20",X"35",X"C0",X"21",
		X"98",X"20",X"7E",X"D3",X"05",X"3A",X"82",X"20",X"A7",X"CA",X"89",X"17",X"2B",X"7E",X"2B",X"77",
		X"2B",X"36",X"01",X"3E",X"04",X"32",X"9B",X"20",X"C9",X"3A",X"98",X"20",X"E6",X"30",X"D3",X"05",
		X"C9",X"3A",X"95",X"20",X"A7",X"CA",X"C6",X"17",X"21",X"F3",X"19",X"11",X"03",X"1A",X"3A",X"82",
		X"20",X"BE",X"D2",X"AA",X"17",X"23",X"13",X"C3",X"A1",X"17",X"1A",X"32",X"97",X"20",X"21",X"98",
		X"20",X"7E",X"E6",X"30",X"47",X"7E",X"E6",X"0F",X"07",X"FE",X"10",X"C2",X"C0",X"17",X"3E",X"01",
		X"B0",X"77",X"AF",X"32",X"95",X"20",X"21",X"99",X"20",X"35",X"C0",X"06",X"EF",X"C3",X"BE",X"19",
		X"3A",X"67",X"20",X"0F",X"D2",X"DA",X"17",X"DB",X"01",X"C9",X"DB",X"02",X"C9",X"DB",X"02",X"E6",
		X"04",X"C8",X"3A",X"9A",X"20",X"A7",X"C0",X"31",X"00",X"24",X"06",X"04",X"CD",X"C5",X"09",X"05",
		X"C2",X"EC",X"17",X"3E",X"01",X"32",X"9A",X"20",X"CD",X"BA",X"19",X"FB",X"11",X"BC",X"1C",X"21");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
