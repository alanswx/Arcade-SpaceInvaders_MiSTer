//============================================================================
//  Arcade: Space Invaders
//
//  Port to MiSTer Dave Wood (oldgit)
//  April 2019 
//
//  This program is free software; you can redistribute it and/or modify it
//  under the terms of the GNU General Public License as published by the Free
//  Software Foundation; either version 2 of the License, or (at your option)
//  any later version.
//
//  This program is distributed in the hope that it will be useful, but WITHOUT
//  ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
//  FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License for
//  more details.
//
//  You should have received a copy of the GNU General Public License along
//  with this program; if not, write to the Free Software Foundation, Inc.,
//  51 Franklin Street, Fifth Floor, Boston, MA 02110-1301 USA.
//============================================================================
module emu
(
	//Master input clock
	input         CLK_50M,

	//Async reset from top-level module.
	//Can be used as initial reset.
	input         RESET,

	//Must be passed to hps_io module
	inout  [45:0] HPS_BUS,

	//Base video clock. Usually equals to CLK_SYS.
	output        VGA_CLK,

	//Multiple resolutions are supported using different VGA_CE rates.
	//Must be based on CLK_VIDEO
	output        VGA_CE,

	output  [7:0] VGA_R,
	output  [7:0] VGA_G,
	output  [7:0] VGA_B,
	output        VGA_HS,
	output        VGA_VS,
	output        VGA_DE,    // = ~(VBlank | HBlank)
	output        VGA_F1,

	//Base video clock. Usually equals to CLK_SYS.
	output        HDMI_CLK,

	//Multiple resolutions are supported using different HDMI_CE rates.
	//Must be based on CLK_VIDEO
	output        HDMI_CE,

	output  [7:0] HDMI_R,
	output  [7:0] HDMI_G,
	output  [7:0] HDMI_B,
	output        HDMI_HS,
	output        HDMI_VS,
	output        HDMI_DE,   // = ~(VBlank | HBlank)
	output  [1:0] HDMI_SL,   // scanlines fx

	//Video aspect ratio for HDMI. Most retro systems have ratio 4:3.
	output  [7:0] HDMI_ARX,
	output  [7:0] HDMI_ARY,

	output        LED_USER,  // 1 - ON, 0 - OFF.

	// b[1]: 0 - LED status is system status OR'd with b[0]
	//       1 - LED status is controled solely by b[0]
	// hint: supply 2'b00 to let the system control the LED.
	output  [1:0] LED_POWER,
	output  [1:0] LED_DISK,

	output [15:0] AUDIO_L,
	output [15:0] AUDIO_R,
	output        AUDIO_S,    // 1 - signed audio samples, 0 - unsigned

	//SDRAM interface with lower latency
	output        SDRAM_CLK,
	output        SDRAM_CKE,
	output [12:0] SDRAM_A,
	output  [1:0] SDRAM_BA,
	inout  [15:0] SDRAM_DQ,
	output        SDRAM_DQML,
	output        SDRAM_DQMH,
	output        SDRAM_nCS,
	output        SDRAM_nCAS,
	output        SDRAM_nRAS,
	output        SDRAM_nWE,  
	
	
		// Open-drain User port.
	// 0 - D+/RX
	// 1 - D-/TX
	// 2..6 - USR2..USR6
	// Set USER_OUT to 1 to read from USER_IN.
	input   [6:0] USER_IN,
	output  [6:0] USER_OUT

);

assign VGA_F1    = 0;
assign USER_OUT  = '1;
assign LED_USER  = ioctl_download;
assign LED_DISK  = 0;
assign LED_POWER = 0;

assign HDMI_ARX = status[1] ? 8'd16 : (status[2] | landscape) ? 8'd4 : 8'd3;
assign HDMI_ARY = status[1] ? 8'd9  : (status[2] | landscape) ? 8'd3 : 8'd4;



`include "build_id.v" 
localparam CONF_STR = {
	"A.INVADERS;;",
	"-;",
	"H0O1,Aspect Ratio,Original,Wide;", 
	"H1H0O2,Orientation,Vert,Horz;",
	"O35,Scandoubler Fx,None,HQ2x,CRT 25%,CRT 50%,CRT 75%;",  
	"-;",
	"DIP;",
	"-;",
	"O8,Overlay,On,Off;",
	"O9,Overlay Test,Off,On;",
	"OA,Background Graphic,On,Off;",
	"-;",
	"H2OBC,Gun Control,Joy1,Joy2,Mouse,Disabled;",
	"H3ODE,Crosshair,Small,Medium,Big,None;",
	"-;",
	"R0,Reset;",
	"J1,Fire 1,Fire 2,Fire 3,Fire 4,Start 1P,Start 2P,Coin;",
	"V,v",`BUILD_DATE
};

////////////////////   CLOCKS   ///////////////////

wire clk_80,clk_40, clk_10;
wire clk_mem = clk_80;
wire clk_sys = clk_10;
wire pll_locked;

pll pll
(
	.refclk(CLK_50M),
	.rst(0),
	.outclk_0(clk_40),
	.outclk_1(clk_10),
	.outclk_2(clk_80),
	.locked(pll_locked)

);


///////////////////////////////////////////////////

wire [31:0] status;
wire  [1:0] buttons;
wire        forced_scandoubler;
wire        direct_video;

wire        ioctl_download;
wire        ioctl_wr;
wire [24:0] ioctl_addr;
wire  [7:0] ioctl_dout;
wire  [7:0] ioctl_index;

reg	[7:0] machine_info;



wire [10:0] ps2_key;
wire [24:0] ps2_mouse;

wire [15:0] joy1, joy2, joy3, joy4;
wire [15:0] joya, joya2;

wire [21:0] gamma_bus;

wire [15:0] sdram_sz;

hps_io #(.STRLEN($size(CONF_STR)>>3)) hps_io
(
   .clk_sys(clk_sys),
   .HPS_BUS(HPS_BUS),

   .conf_str(CONF_STR),

   .buttons(buttons),
   .status(status),
   .status_menumask({&gun_mode|!gun_game,!gun_game,landscape,direct_video}),
   .forced_scandoubler(forced_scandoubler),
   .gamma_bus(gamma_bus),
   .direct_video(direct_video),

   .ioctl_download(ioctl_download),
   .ioctl_wr(ioctl_wr),
   .ioctl_addr(ioctl_addr),
   .ioctl_dout(ioctl_dout),
   .ioctl_index(ioctl_index),

   .sdram_sz(sdram_sz),

	
   .joystick_0(joy1),
   .joystick_1(joy2),
   .joystick_2(joy3),
   .joystick_3(joy4),
   .joystick_analog_0(joya),
   .joystick_analog_1(joya2),
   .ps2_key(ps2_key),
	.ps2_mouse(ps2_mouse)
);

wire       pressed = ps2_key[9];
wire [8:0] code    = ps2_key[8:0];
always @(posedge clk_sys) begin
	reg old_state;
	old_state <= ps2_key[10];
	
	if(old_state != ps2_key[10]) begin
		casex(code)
			'h75: btn_up            <= pressed; // up
			'h72: btn_down          <= pressed; // down
			'h6B: btn_left          <= pressed; // left
			'h74: btn_right         <= pressed; // right
			'h76: btn_coin1         <= pressed; // ESC
			'h05: btn_start1        <= pressed; // F1
			'h06: btn_start2        <= pressed; // F2
			'h14: btn_fireA         <= pressed; // lctrl
			'h11: btn_fireB         <= pressed; // lalt
			'h29: btn_fireC         <= pressed; // Space
			'h12: btn_fireD         <= pressed; // l-shift

			// JPAC/IPAC/MAME Style Codes
			'h16: btn_start1        <= pressed; // 1
			'h1E: btn_start2        <= pressed; // 2
                        'h26: btn_start3        <= pressed; // 3
			'h25: btn_start4        <= pressed; // 4

			'h2E: btn_coin1         <= pressed; // 5
			'h36: btn_coin2         <= pressed; // 6
			'h2D: btn_up2           <= pressed; // R
			'h2B: btn_down2         <= pressed; // F
			'h23: btn_left2         <= pressed; // D
			'h34: btn_right2        <= pressed; // G
			'h1C: btn_fire2A        <= pressed; // A
			'h1B: btn_fire2B        <= pressed; // S
			'h21: btn_fire2C        <= pressed; // Q
			'h1D: btn_fire2D        <= pressed; // W
		endcase
	end
end


reg btn_left   = 0;
reg btn_right  = 0;
reg btn_down   = 0;
reg btn_up     = 0;
reg btn_fireA  = 0;
reg btn_fireB  = 0;
reg btn_fireC  = 0;
reg btn_fireD  = 0;
reg btn_coin1  = 0;
reg btn_coin2  = 0;
reg btn_start1 = 0;
reg btn_start2 = 0;
reg btn_start3 = 0;
reg btn_start4 = 0;
reg btn_up2    = 0;
reg btn_down2  = 0;
reg btn_left2  = 0;
reg btn_right2 = 0;
reg btn_fire2A = 0;
reg btn_fire2B = 0;
reg btn_fire2C = 0;
reg btn_fire2D = 0;

wire m_start1  = btn_start1 | joy[8];
wire m_start2  = btn_start2 | joy[9];
wire m_coin1   = btn_coin1  | btn_coin2 | joy[10];

wire m_right1  = btn_right  | joy1[0];
wire m_left1   = btn_left   | joy1[1];
wire m_down1   = btn_down   | joy1[2];
wire m_up1     = btn_up     | joy1[3];
wire m_fire1a  = btn_fireA  | joy1[4] | ps2_mouse[0];
wire m_fire1b  = btn_fireB  | joy1[5] | ps2_mouse[1];
wire m_fire1c  = btn_fireC  | joy1[6] | ps2_mouse[2];
wire m_fire1d  = btn_fireD  | joy1[7];

wire m_right2  = btn_right2 | joy2[0];
wire m_left2   = btn_left2  | joy2[1];
wire m_down2   = btn_down2  | joy2[2];
wire m_up2     = btn_up2    | joy2[3];
wire m_fire2a  = btn_fire2A | joy2[4];
wire m_fire2b  = btn_fire2B | joy2[5];
wire m_fire2c  = btn_fire2C | joy2[6];
wire m_fire2d  = btn_fire2D | joy2[7];

wire m_right   = m_right1 | m_right2;
wire m_left    = m_left1  | m_left2; 
wire m_down    = m_down1  | m_down2; 
wire m_up      = m_up1    | m_up2;   
wire m_fire_a  = m_fire1a | m_fire2a;
wire m_fire_b  = m_fire1b | m_fire2b;
wire m_fire_c  = m_fire1c | m_fire2c;
wire m_fire_d  = m_fire1d | m_fire2d;

wire m_coin3   = joy3[10];
wire m_start3  = joy3[8] | btn_start3;
wire m_left3   = joy3[1];
wire m_right3  = joy3[0];
wire m_up3     = joy3[3];
wire m_down3   = joy3[2];
/*
wire m_fire3a  = joy3[4];
wire m_fire3b  = joy3[5];
wire m_fire3c  = joy3[6];
wire m_fire3d  = joy3[7];
*/

wire m_coin4   = joy4[10];
wire m_start4  = joy4[8] | btn_start4;
wire m_left4   = joy4[1];
wire m_right4  = joy4[0];
wire m_up4     = joy4[3];
wire m_down4   = joy4[2];
/*
wire m_fire4a  = joy4[4];
wire m_fire4b  = joy4[5];
wire m_fire4c  = joy4[6];
wire m_fire4d  = joy4[7];
*/


wire [2:0] ms_col;
wire [2:0] bs_col;
wire [2:0] sh_col;
wire [2:0] sc1_col;
wire [2:0] sc2_col;
wire [2:0] mn_col;

wire [15:0] joy = joy1 | joy2;


///////////////////////////////////////////////////////////////////


wire hblank;
wire vblank;
//wire hs, vs;
wire r,g,b;
//wire no_rotate = 1'b1;//status[2] | direct_video | landscape;
wire no_rotate = status[2] | direct_video | landscape;
reg ce_pix;
always @(posedge clk_40) begin
        reg [2:0] div;

        div <= div + 1'd1;
	ce_pix <= div == 0;
end

wire fg = |{rr,gg,bb};

wire [7:0]rr = {8{r}};
wire [7:0]gg = {8{g}};
wire [7:0]bb = {8{b}};

// if graphics are turned off, just use the pixels. Otherwise if the
// background is in effect - use it
wire [23:0] rgbdata  = (gun_target & (~&gun_mode & gun_game)) ? {8'd255, 16'd0} : status[10]? {rr,gg,bb}  : (fg && !bg_a) ? {rr,gg,bb} : {bg_r,bg_g,bg_b};



//arcade_video #(260,224,6) arcade_video
arcade_video #(260,224,24) arcade_video
(
   .*,

   .clk_video(clk_40),

  // .RGB_in({r,r,g,g,b,b}),
   //.RGB_in((fg && !bg_a) ? {rr,gg,bb} : {bg_r,bg_g,bg_b}),
   .RGB_in(rgbdata),
   //.RGB_in({bg_r,bg_g,bg_b}),
   //.RGB_in(status[10]?  {bg_r,bg_g,bg_b}:{rr,gg,bb}  ),

   .HBlank(hblank),
   .VBlank(vblank),
   .HSync(HSync),
   .VSync(VSync),

   .rotate_ccw(ccw),
   .fx(status[5:3])

);


wire [7:0] audio;
wire [7:0] inv_audio_data;
wire [7:0] zap_audio_data;

assign AUDIO_L = (mod==mod_280zap)? {zap_audio_data,zap_audio_data}:{inv_audio_data,inv_audio_data};

//assign AUDIO_L = {audio, audio};
assign AUDIO_R = AUDIO_L;
assign AUDIO_S = 0;
wire reset;
assign reset = (RESET | status[0] | buttons[1] | ioctl_download);

wire [7:0] GDB0;
wire [7:0] GDB1;
wire [7:0] GDB2;
wire [7:0] GDB3;
wire [7:0] GDB4;
wire [7:0] GDB5;
wire [7:0] GDB6;


localparam mod_spaceinvaders = 0;
localparam mod_shuffleboard  = 1;
localparam mod_vortex        = 2;
localparam mod_280zap        = 3;
localparam mod_blueshark     = 4;
localparam mod_boothill      = 5;
localparam mod_lunarrescue   = 6;
localparam mod_ozmawars      = 7;
localparam mod_spacelaser    = 8;
localparam mod_spacewalk     = 9;
localparam mod_spaceinvaderscv = 10;
localparam mod_unknown1      = 11;
localparam mod_unknown2      = 12;
localparam mod_spaceinvadersii = 13;
localparam mod_amazingmaze   = 14;
localparam mod_attackforce   = 15;
localparam mod_ballbomb      = 16;
localparam mod_bowler        = 17;
localparam mod_checkmate     = 18;
localparam mod_clowns        = 19;
localparam mod_cosmo         = 20;
localparam mod_dogpatch      = 21;
localparam mod_doubleplay    = 22;
localparam mod_guidedmissle  = 23;
localparam mod_claybust      = 24;
localparam mod_gunfight      = 25;
localparam mod_indianbattle  = 26;
localparam mod_lupin         = 27;
localparam mod_m4            = 28;
localparam mod_phantom       = 29;
localparam mod_polaris       = 30;
localparam mod_desertgun     = 31;
localparam mod_lagunaracer   = 32;
localparam mod_seawolf       = 33;
localparam mod_yosakdon      = 34;
localparam mod_spacechaser   = 35;
localparam mod_steelworker   = 36;


reg [7:0] mod = 0;
always @(posedge clk_sys) if (ioctl_wr & (ioctl_index==1)) mod <= ioctl_dout;

 
wire [9:0] center_joystick_y   =  8'd127 + joya[15:8];
//wire [9:0] positive_joystick_y   =  joya[15] ? 8'd128+ $signed(joya[15:8]) : 10'b0;
wire [7:0] positive_joystick_y   =  joya[15] ? ~joya[15:8] : 10'b0;
wire [7:0] positive_joystick_y_2   =  joya2[15] ? ~joya2[15:8] : 10'b0;
wire   [3:0] zap_throttle = positive_joystick_y[6:3] ;

/* controls for blue shark */
wire [7:0] bluerange = { 1'b0, gun_x[7:1]+8'd8 };
reg [7:0] blue_shark_x;

always @(posedge clk_sys) 
begin
   if (bluerange > 9'h082)
	   blue_shark_x=8'h82;
   else
	   blue_shark_x=bluerange[7:0];
end

/* controls for claybust */
wire [15:0] gun_x_16 = gun_x;
wire [15:0] gun_y_16 = gun_y + 8'h20;
wire [15:0] claybust_gun_pos = (((gun_x_16 >> 3) | (gun_y_16 << 5)) + 2);
reg [7:0] claybust_gun_pos_lo;
reg [7:0] claybust_gun_pos_hi;
reg [19:0] claybust_gun_on;
reg claybust_old_fire;
always @(posedge clk_10) begin
	claybust_gun_pos_lo <= claybust_gun_pos & 8'hff;
	claybust_gun_pos_hi <= claybust_gun_pos >> 8;
	claybust_old_fire <= m_fire1a;
	if (~claybust_old_fire & m_fire1a) claybust_gun_on <= 20'hfffff; // arbitrary
	else if (claybust_gun_on) claybust_gun_on <= claybust_gun_on - 1;
end

/* controls for desert gun */
reg [7:0] desert_gun_x;
reg [7:0] desert_gun_y;
reg desert_gun_select;

always @(posedge clk_sys) 
begin
	desert_gun_x <= (gun_x[7:0]>>1)+8'h10;
	desert_gun_y <= (gun_y[7:0]>>1)+8'h10;
	if (Trigger_AudioDeviceP2) desert_gun_select <= SoundCtrl5[3];
end

/* controls for clown */
reg [7:0] clown_y = 128;
reg [5:0] clown_timer= 0;
reg vsync_r;
//always @(posedge m_right or posedge m_left ) begin
always @(posedge clk_sys) 
begin
    vsync_r          <= VSync;
    if (vsync_r ==0 && VSync== 1) 
    begin
       //if (clown_timer > 1) begin
        if (m_right && clown_y < 255)
            clown_y <= clown_y +1;
        else if (m_left && clown_y > 0)
            clown_y <= clown_y -1;
       clown_timer <= clown_timer +1;
       //end
       //else
	//     clown_timer <= clown_timer +1;
    end
end

/* controls for dogpatch */
/* dogpatch has some weird non incremental thing going on*/
/*0x07, 0x06, 0x04, 0x05, 0x01, 0x00, 0x02*/
/* gunfight */
/*0x06, 0x02, 0x00, 0x04, 0x05, 0x01, 0x03*/
reg [2:0] dogpatch_y_count= 0;
reg [2:0] dogpatch_y_2_count= 0;
reg [2:0] gunfight_y_count= 0;
reg [2:0] gunfight_y_count_2= 0;
wire [2:0] dogpatch_y;
wire [2:0] dogpatch_y_2;
wire [2:0] gunfight_y;
wire [2:0] gunfight_y_2;
reg [5:0] dogpatch_timer= 0;
always @(posedge clk_sys) 
begin
    if (vsync_r ==0 && VSync== 1) 
    begin
	if (dogpatch_timer == 8'd5) 
	begin
          if (m_up&& dogpatch_y_count< 7)
            dogpatch_y_count<= dogpatch_y_count+1;
          else if (m_down&& dogpatch_y_count > 0)
            dogpatch_y_count<= dogpatch_y_count-1;

          if (m_up2&& dogpatch_y_2_count< 7)
            dogpatch_y_2_count<= dogpatch_y_2_count+1;
          else if (m_down2&& dogpatch_y_2_count > 0)
            dogpatch_y_2_count<= dogpatch_y_2_count-1;

          if (m_fire1b&& gunfight_y_count< 7)
            gunfight_y_count<= gunfight_y_count+1;
          else if (m_fire1c&& gunfight_y_count > 0)
            gunfight_y_count<= gunfight_y_count-1;

          if (m_fire2b&& gunfight_y_count_2< 7)
            gunfight_y_count_2<= gunfight_y_count_2+1;
          else if (m_fire2c&& gunfight_y_count_2 > 0)
            gunfight_y_count_2<= gunfight_y_count_2-1;


          dogpatch_timer <= 0;
        end
	else 
	begin
          dogpatch_timer <= dogpatch_timer +1;
	end
        case (dogpatch_y_count) 
		3'b000: dogpatch_y <= 3'h7;
		3'b001: dogpatch_y <= 3'h6;
		3'b010: dogpatch_y <= 3'h4;
		3'b011: dogpatch_y <= 3'h5;
		3'b100: dogpatch_y <= 3'h1;
		3'b101: dogpatch_y <= 3'h0;
		3'b110: dogpatch_y <= 3'h2;
		3'b111: dogpatch_y <= 3'h2; // ?
	endcase
        case (dogpatch_y_2_count) 
		3'b000: dogpatch_y_2 <= 3'h7;
		3'b001: dogpatch_y_2 <= 3'h6;
		3'b010: dogpatch_y_2 <= 3'h4;
		3'b011: dogpatch_y_2 <= 3'h5;
		3'b100: dogpatch_y_2 <= 3'h1;
		3'b101: dogpatch_y_2 <= 3'h0;
		3'b110: dogpatch_y_2 <= 3'h2;
		3'b111: dogpatch_y_2 <= 3'h2; // ?
	endcase
        case (gunfight_y_count) 
		3'b000: gunfight_y <= 3'h6;
		3'b001: gunfight_y <= 3'h2;
		3'b010: gunfight_y <= 3'h0;
		3'b011: gunfight_y <= 3'h4;
		3'b100: gunfight_y <= 3'h5;
		3'b101: gunfight_y <= 3'h1;
		3'b110: gunfight_y <= 3'h3;
		3'b111: gunfight_y <= 3'h3; //?
	endcase
        case (gunfight_y_count_2) 
		3'b000: gunfight_y_2 <= 3'h6;
		3'b001: gunfight_y_2 <= 3'h2;
		3'b010: gunfight_y_2 <= 3'h0;
		3'b011: gunfight_y_2 <= 3'h4;
		3'b100: gunfight_y_2 <= 3'h5;
		3'b101: gunfight_y_2 <= 3'h1;
		3'b110: gunfight_y_2 <= 3'h3;
		3'b111: gunfight_y_2 <= 3'h3; //?
	endcase
    end
end

/* controls for seawolf */
wire [7:0] seawolf_shifted_x = gun_x[7:0]>>3;
reg [4:0] seawolf_position;

always @(posedge clk_sys) 
begin
   case (seawolf_shifted_x[4:0]) 
      5'b00000: seawolf_position <= ~5'h1e; // clamp
      5'b00001: seawolf_position <= ~5'h1e;
      5'b00010: seawolf_position <= ~5'h1c;
      5'b00011: seawolf_position <= ~5'h1d;
      5'b00100: seawolf_position <= ~5'h19;
      5'b00101: seawolf_position <= ~5'h18;
      5'b00110: seawolf_position <= ~5'h1a;
      5'b00111: seawolf_position <= ~5'h1b;
      5'b01000: seawolf_position <= ~5'h13;
      5'b01001: seawolf_position <= ~5'h12;
      5'b01010: seawolf_position <= ~5'h10;
      5'b01011: seawolf_position <= ~5'h11;
      5'b01100: seawolf_position <= ~5'h15;
      5'b01101: seawolf_position <= ~5'h14;
      5'b01110: seawolf_position <= ~5'h16;
      5'b01111: seawolf_position <= ~5'h17;
      5'b10000: seawolf_position <= ~5'h07;
      5'b10001: seawolf_position <= ~5'h06;
      5'b10010: seawolf_position <= ~5'h04;
      5'b10011: seawolf_position <= ~5'h05;
      5'b10100: seawolf_position <= ~5'h01;
      5'b10101: seawolf_position <= ~5'h00;
      5'b10110: seawolf_position <= ~5'h02;
      5'b10111: seawolf_position <= ~5'h03;
      5'b11000: seawolf_position <= ~5'h0b;
      5'b11001: seawolf_position <= ~5'h0a;
      5'b11010: seawolf_position <= ~5'h08;
      5'b11011: seawolf_position <= ~5'h09;
      5'b11100: seawolf_position <= ~5'h0d;
      5'b11101: seawolf_position <= ~5'h0c;
      5'b11110: seawolf_position <= ~5'h0e;
      5'b11111: seawolf_position <= ~5'h0e; // clamp
   endcase
end

reg fire_toggle = 0;
always @(posedge m_fire_a) fire_toggle <= ~fire_toggle;

reg [7:0] sw[8];
always @(posedge clk_sys) if (ioctl_wr && (ioctl_index==254) && !ioctl_addr[24:3]) sw[ioctl_addr[2:0]] <= ioctl_dout;

reg landscape;
reg ccw;
reg color_rom_enabled;

wire WDEnabled;
wire Trigger_ShiftCount;
wire Trigger_ShiftData;
wire Trigger_AudioDeviceP1;
wire Trigger_AudioDeviceP2;
wire Trigger_WatchDogReset;
wire [7:0] PortWr;
wire [7:0] S;
wire [7:0] SR= { S[0], S[1], S[2], S[3], S[4], S[5], S[6], S[7]} ;
wire ShiftReverse;

always @(*) begin

        gun_game <= 0;
        landscape <= 1;
        ccw<=0;
        color_rom_enabled<=0;
	WDEnabled <= 1'b1;
        GDB0 <= 8'hFF;
        GDB1 <= 8'hFF;
        GDB2 <= 8'hFF;
        GDB3 <= S;

        // space invaders default PortWr mapping
        Trigger_ShiftCount     <= PortWr[2];
        Trigger_AudioDeviceP1  <= PortWr[3];
        Trigger_ShiftData      <= PortWr[4];
        Trigger_AudioDeviceP2  <= PortWr[5];
        Trigger_WatchDogReset  <= PortWr[6];


        case (mod) 
        mod_spaceinvaders:
        begin
          landscape<=0;
          ccw<=1;

          GDB0 <= sw[0] | { 1'b1, m_right,m_left,m_fire_a,1'b1,1'b1, 1'b1,1'b1};
          GDB1 <= sw[1] | { 1'b1, m_right,m_left,m_fire_a,1'b1,m_start1, m_start2, m_coin1 };
          GDB2 <= sw[2] | { 1'b1, m_right,m_left,m_fire_a,1'b0,1'b0, 1'b1, 1'b1 };
        end
        mod_shuffleboard:
        begin
          landscape<=0;
          ccw<=0;
          GDB1 <= S;
	  // IN0
          GDB2 <= sw[1] | ~{ 1'b0, m_right,m_left,m_fire_a,1'b0,m_start1, m_start2, m_coin1 };
          GDB3 <= SR;
	  // IN1
	  // GB4 <=
	  // IN2 // trackball Y
	  // GB5 <=
	  // IN3 // trackball X
	  // GB6 <=
	  // 4,5,6 ???
          Trigger_ShiftCount     <= PortWr[1];
          Trigger_AudioDeviceP1  <= PortWr[5];
          Trigger_ShiftData      <= PortWr[2];
          Trigger_AudioDeviceP2  <= PortWr[6];
          Trigger_WatchDogReset  <= PortWr[4];
        end
        mod_vortex:
        begin
          //GDB0 -- all FF
          //
          landscape<=0;
          ccw<=1;
	  // IN2 -- settings
          GDB0 <= sw[2] | { 1'b0, m_right2,m_left2,m_fire2a,1'b0,1'b0, 1'b0, 1'b0};
          GDB1 <= S;
	  // IN0
	  //GDB2 <= sw[1] | { 1'b1, m_right1,m_left1,m_fire1a,1'b1,m_start1, m_start2, ~m_coin1 };
	  //GDB2 <= sw[1] | { 1'b1, m_right1,m_left1,m_fire1a,1'b1,m_start1, m_start2, ~m_coin1 };
          GDB2 <= 8'h00;
	  // IN1
          GDB3 <= sw[1] | { 1'b0, m_right2,m_left2,m_fire2a,1'b0,m_start1, m_start2, ~m_coin1 };
	  
          Trigger_ShiftCount     <= PortWr[0];
          Trigger_AudioDeviceP1  <= PortWr[1];
          Trigger_ShiftData      <= PortWr[6];
          Trigger_AudioDeviceP2  <= PortWr[7];
          Trigger_WatchDogReset  <= PortWr[4];
        end
        mod_lagunaracer:
	begin
 	  landscape<=0;
	   GDB0 <= sw[0] | { ~m_start1, ~m_coin1, 1'b1, fire_toggle, zap_throttle};
           //GDB1 <= sw[1] | { 1'b0, 1'b1, 1'b1,1'b1,1'b1,1'b1, 1'b1, 1'b1 };
           GDB1 <= 8'd127-joya[7:0];
           GDB2 <= sw[2] | { 1'b0, 1'b0, 1'b0,1'b0,1'b0,1'b0, 1'b0, 1'b0 };
	  // IN0
          //GDB0 <= sw[0] | { m_start1, m_coin1,1'b1,m_fire_a,1'b1,1'b0, 1'b0,1'b0};
	  // IN1
          //GDB1 <= sw[1] | { 1'b0, 1'b1,1'b1,1'b1,1'b1,1'b1, 1'b1, 1'b1 };
	  // IN2
          //GDB2 <= sw[2] | { 1'b1, 1'b1,1'b0,1'b0,1'b0,1'b0, 1'b0, 1'b0 };
          Trigger_ShiftCount     <= PortWr[4];
          Trigger_AudioDeviceP1  <= PortWr[2];
          Trigger_ShiftData      <= PortWr[3];
          Trigger_AudioDeviceP2  <= PortWr[5];
          Trigger_WatchDogReset  <= PortWr[7];
        end
	mod_280zap:
	begin
 	  landscape<=1;
	   //GDB0 <= sw[0] | { ~m_start1, ~m_coin1, 1'b1, m_fire_a, m_fire_b,1'b0,1'b0,1'b0/*(joya[11:8]*/};
	   GDB0 <= sw[0] | { ~m_start1, ~m_coin1, 1'b1, fire_toggle, zap_throttle};
           //GDB1 <= sw[1] | { 1'b0, 1'b1, 1'b1,1'b1,1'b1,1'b1, 1'b1, 1'b1 };
           GDB1 <= 8'd127-joya[7:0];
           GDB2 <= sw[2] | { 1'b0, 1'b0, 1'b0,1'b0,1'b0,1'b0, 1'b0, 1'b0 };
	  // IN0
          //GDB0 <= sw[0] | { m_start1, m_coin1,1'b1,m_fire_a,1'b1,1'b0, 1'b0,1'b0};
	  // IN1
          //GDB1 <= sw[1] | { 1'b0, 1'b1,1'b1,1'b1,1'b1,1'b1, 1'b1, 1'b1 };
	  // IN2
          //GDB2 <= sw[2] | { 1'b1, 1'b1,1'b0,1'b0,1'b0,1'b0, 1'b0, 1'b0 };
          Trigger_ShiftCount     <= PortWr[4];
          Trigger_AudioDeviceP1  <= PortWr[2];
          Trigger_ShiftData      <= PortWr[3];
          Trigger_AudioDeviceP2  <= PortWr[5];
          Trigger_WatchDogReset  <= PortWr[7];

	end

        mod_blueshark:
        begin
		    gun_game <= 1;
          GDB0 <= SR;
	  // IN0
          //GDB1 <= 8'd127-joya[7:0];
          //GDB1 <= { 8'b01000010};
        //  GDB1 <= { 8'd63 + joya[7:1]};

          //GDB1 <= (blue_control[8:1]+8'd8) ;
          GDB1 <= blue_shark_x;
	  // IN1
          GDB2 <= sw[2] | { 1'b0, 1'b0,1'b0,1'b1,1'b1,1'b1,m_coin1 ,~m_fire_a};
          Trigger_ShiftCount     <= PortWr[1];
          Trigger_AudioDeviceP1  <= PortWr[3];
          Trigger_ShiftData      <= PortWr[2];
          Trigger_WatchDogReset  <= PortWr[4];
        end
        mod_boothill:
        begin 
          // IN0
          GDB0 <= sw[0] | { m_fire1a, 1'b0,1'b1,1'b0,m_right1,m_left1,m_down1,m_up1};
          // IN1
          GDB1 <= sw[1] | { m_fire2a, 1'b0,1'b1,1'b0,m_right2,m_left2,m_down2,m_up2};
          // IN2
          GDB2 <= sw[2] | { m_start1, m_coin1,m_start1,1'b0,1'b1,1'b1, 1'b0, 1'b1 };
          Trigger_ShiftCount     <= PortWr[1]; // IS THIS WEIRD?
          Trigger_AudioDeviceP1  <= PortWr[3];
          Trigger_ShiftData      <= PortWr[2];
          Trigger_WatchDogReset  <= PortWr[4];
          //<= PortWr[5]; // tone_generator_low_w
          //<= PortWr[6]; // tone_generator_hi_w
	  GDB3 <= ShiftReverse ? SR: S;

        end
        mod_lunarrescue:
        begin
          landscape<=0;
          color_rom_enabled<=1;
          ccw<=1;
	  WDEnabled <= 1'b0;
          //GDB0 <= sw[0] | { 1'b1, m_right,m_left,m_fire_a,1'b1,1'b0, 1'b0,1'b0};
          //GDB1 <= sw[1] | { 1'b1, m_right,m_left,m_fire_a,1'b1,m_start1, m_start2, m_coin1 };
          //GDB2 <= sw[2] | { 1'b1, m_right,m_left,m_fire_a,1'b0,1'b0, 1'b1, 1'b1 };
          GDB0 <= sw[0] | { 1'b1, 1'b0,1'b0,1'b0,1'b0,1'b1, 1'b0,1'b0};
          //GDB0 <= sw[0] | { 1'b0, 1'b0, 1'b0, m_right,m_left,m_fire_a,1'b1,1'b1, 1'b1,1'b1};
          GDB1 <= sw[1] | { 1'b1, m_right,m_left,m_fire_a,1'b0,m_start1, m_start2, ~m_coin1 };
          GDB2 <= sw[2] | { 1'b1, m_right,m_left,m_fire_a,1'b0,1'b0, 1'b1, 1'b1 };
        end
        mod_ozmawars:
        begin
            landscape<=0;
            ccw<=1;
            color_rom_enabled<=1;
         // GDB0 <= sw[0] | ~{ 1'b0, m_right,m_left,m_fire_a,1'b0,1'b1, 1'b1,1'b1};
            GDB1 <= sw[1] | { 1'b1, m_right,m_left,m_fire_a,1'b0,m_start1, m_start2, ~m_coin1 };
            GDB2 <= sw[2] | { m_start1, m_coin1,m_start2,1'b0,1'b0,1'b0, 1'b0, 1'b0 };
          end
        mod_spacelaser:
        begin
            landscape<=0;
            ccw<=1;
            color_rom_enabled<=1;
        // GDB0 <= sw[0] | ~{ 1'b0, m_right,m_left,m_fire_a,1'b0,1'b1, 1'b1,1'b1};
            GDB1 <= sw[1] | { 1'b1, m_right,m_left,m_fire_a,1'b1,m_start1, m_start2, m_coin1 };
            GDB2 <= sw[2] | { 1'b1, m_right,m_left,m_fire_a,1'b0,1'b0, 1'b0, 1'b0 };
		  end
        mod_spacewalk:
        begin
	     WDEnabled <= 1'b0;
             GDB0 <= clown_y;
             GDB1 <= sw[1] | { 1'b1,~m_coin1,~m_start1,~m_start2,1'b1,1'b1,1'b1,1'b1};
             GDB2 <= sw[2];
             Trigger_ShiftCount     <= PortWr[1];
             Trigger_AudioDeviceP1  <= PortWr[3];
             Trigger_ShiftData      <= PortWr[2];
             Trigger_AudioDeviceP2  <= PortWr[6];
             Trigger_WatchDogReset  <= PortWr[7];
             //<= PortWr[5]; // tone_generator_low_w
             //<= PortWr[6]; // tone_generator_hi_w
        end
        mod_spaceinvaderscv:
        begin
            landscape<=0;
            ccw<=1;
            color_rom_enabled<=1;
            GDB0 <= sw[0] | { 1'b0, 1'b0,1'b0,1'b0,1'b0,1'b0, 1'b0,1'b0};
            GDB1 <= sw[1] | { 1'b1, m_right,m_left,m_fire_a,1'b1,m_start1, m_start2, m_coin1 };
            GDB2 <= sw[2] | { 1'b1, m_right,m_left,m_fire_a,1'b0,1'b0, 1'b0, 1'b0 };
        end
        mod_unknown1:
        begin
        GDB0 <= 8'hFF;
        GDB1 <= 8'hFF;
        GDB2 <= 8'hFF;
        end
        mod_unknown2:
        begin
        GDB0 <= 8'h00;
        GDB1 <= 8'h00;
        GDB2 <= 8'h00;
        end
        mod_spaceinvadersii:
        begin
	 landscape<=0;
          ccw<=1;
          color_rom_enabled<=1;
          GDB0 <= sw[0] | { 1'b0, 1'b0,1'b0,1'b0,1'b0,1'b1, 1'b0,1'b0};
          //GDB0 <= sw[0] | { 1'b0, 1'b0, 1'b0, m_right,m_left,m_fire_a,1'b1,1'b1, 1'b1,1'b1};
          GDB1 <= sw[1] | { 1'b1, m_right,m_left,m_fire_a,1'b0,m_start1, m_start2, ~m_coin1 };
          GDB2 <= sw[2] | { 1'b1, m_right,m_left,m_fire_a,1'b0,1'b0, 1'b1, 1'b1 };
        end
        mod_amazingmaze:
        begin
	     WDEnabled <= 1'b0;
             GDB0 <= sw[0] | { m_up2, m_down2, m_right2, m_left2, m_up1, m_down1, m_right1, m_left1} ;
             GDB1 <= sw[1] | { 1'b0, 1'b0,1'b0,1'b0,m_coin1, 1'b0, m_start2, m_start1};
             GDB2 <= 8'b0;
        end
        mod_attackforce:
	begin
            landscape<=1;
	    WDEnabled <= 1'b0;
            ccw<=1;
            GDB0 <= sw[0] | { ~m_coin1, 1'b1,1'b1,1'b1,1'b1,~m_fire_a, ~m_left,~m_right};
            GDB1 <= 8'b0;
            GDB2 <= 8'b0;
            Trigger_ShiftCount     <= PortWr[7];
            Trigger_AudioDeviceP1  <= PortWr[4];
            Trigger_ShiftData      <= PortWr[3];
            Trigger_AudioDeviceP2  <= PortWr[6];
            Trigger_WatchDogReset  <= PortWr[5];

	end
        mod_ballbomb:
	begin
            landscape<=0;
	    WDEnabled <= 1'b0;
            ccw<=1;
            color_rom_enabled<=1;
            GDB0 <= sw[0] | { 1'b1, m_right,m_left,m_fire_a,1'b0,1'b0, 1'b0, 1'b0 };
            GDB1 <= sw[1] | { 1'b1, m_right,m_left,m_fire_a,1'b1,m_start1, m_start2, m_coin1 };
            GDB2 <= sw[2] | { 1'b0, 1'b0,1'b0,1'b0,1'b0,1'b0, 1'b0,1'b0};
	end
        mod_bowler:
	begin
            landscape<=0;
	// 0 - dips
            GDB0 <= sw[0];
	// 1 - controls
	   GDB1 <= ~S;
            //GDB1 <= sw[1] | { 1'b0,1'b0,1'b0,1'b0,m_fire_b,m_start1, m_fire_a, m_coin1 };
    	// 2, 3 trackball
            GDB2 <= sw[2];
            GDB3 <= ~SR;
             Trigger_ShiftCount     <= PortWr[1];
             //Trigger_AudioDeviceP1  <= PortWr[3];
             Trigger_ShiftData      <= PortWr[2];
             //Trigger_AudioDeviceP2  <= PortWr[6];
             Trigger_WatchDogReset  <= PortWr[4];
             //<= PortWr[5]; // bowler_audio_1_w 
             //<= PortWr[6]; // bowler_audio_2_w
             //<= PortWr[7]; // bowler_lights_1_w
             //<= PortWr[8]; //
             //<= PortWr[9]; //
             //<= PortWr[A]; //
             //<= PortWr[E]; //
             //<= PortWr[F]; //
	end
        mod_checkmate:
	begin
	  WDEnabled <= 1'b0;
          // IN0
          GDB0 <= sw[0] | { m_right2,m_left2,m_down2,m_up2,m_right1,m_left1,m_down1,m_up1};
          GDB1 <= sw[1] | { m_right4,m_left4,m_down4,m_up4,m_right3,m_left3,m_down3,m_up3};
          GDB1 <= sw[1] ;
          GDB2 <= sw[2]; // dips
          GDB3 <= sw[3] | { m_coin1, 1'b0,1'b0,1'b0,m_start4,m_start3,m_start2,m_start1};
          //GDB3 <= sw[3] | { m_coin1, 1'b0,1'b0,1'b0,1'b0,1'b0,m_start2,m_start1};
          //<= PortWr[3]; //  checkmat_io_w
	end
        mod_clowns:
	begin
          //GDB0 -- all FF
          //
          landscape<=1;
	  // IN0
          //GDB0 <= sw[0] | 8'b0;
          //GDB0 <= 8'd127-joya[7:0];
          GDB0 <= clown_y;
          GDB1 <= sw[1] | { 1'b1,~m_coin1,~m_start1,~m_start2,1'b1,1'b1,1'b1,1'b1};
          GDB2 <= sw[2] | { m_up, 1'b0,1'b0,1'b0,1'b0,1'b1, 1'b0,1'b0};
	  
          Trigger_ShiftCount     <= PortWr[1];
          Trigger_AudioDeviceP1  <= PortWr[3];
          Trigger_ShiftData      <= PortWr[2];
          Trigger_AudioDeviceP2  <= PortWr[7];
          Trigger_WatchDogReset  <= PortWr[4];
             //<= PortWr[5]; // tone_generator_low_w
             //<= PortWr[6]; // tone_generator_hi_w
	end
        mod_cosmo:
	begin
            landscape<=0;
            ccw<=0;
            color_rom_enabled<=1;
            GDB0 <= sw[0] | { 1'b0, 1'b0,1'b0,1'b0,1'b0,1'b0, 1'b0,1'b0};
            GDB1 <= sw[1] | { 1'b0, m_right,m_left,m_fire_a,1'b1,m_start1, m_start2, m_coin1 };
            GDB2 <= sw[2] | { 1'b1, m_right,m_left,m_fire_a,1'b0,1'b0, 1'b0, 1'b0 };
        Trigger_ShiftCount     <= 1'b0;
        Trigger_AudioDeviceP1  <= PortWr[3];
        Trigger_ShiftData      <= 1'b0;
        Trigger_AudioDeviceP2  <= PortWr[5];
        Trigger_WatchDogReset  <= PortWr[6];
	end
	mod_dogpatch:
        begin
            landscape<=1;
            ccw<=0;
            color_rom_enabled<=1;
            GDB0 <= sw[0] | { ~m_fire_b, dogpatch_y_2, 1'b1, ~m_start2, ~m_start1, ~m_coin1 };
            GDB1 <= sw[1] | { ~m_fire_a, dogpatch_y, 1'b1, 1'b1, 1'b1 , 1'b1};
            GDB2 <= sw[2];
          Trigger_ShiftCount     <= PortWr[1];
          Trigger_AudioDeviceP1  <= PortWr[3];
          Trigger_ShiftData      <= PortWr[2];
          Trigger_AudioDeviceP2  <= PortWr[7];
          Trigger_WatchDogReset  <= PortWr[4];
             //<= PortWr[5]; // tone_generator_low_w
             //<= PortWr[6]; // tone_generator_hi_w

	end
	mod_doubleplay:
        begin
            landscape<=1;
            ccw<=0;
            color_rom_enabled<=1;
            GDB0 <= sw[0] | { ~m_start1, joya[7:2], ~m_fire_a};
            GDB1 <= sw[1] | { ~m_start2, joya[7:2], ~m_fire_a};
            GDB2 <= sw[2] | { ~m_coin1, 7'b0 };
          Trigger_ShiftCount     <= PortWr[1];
          Trigger_AudioDeviceP1  <= PortWr[3];
          Trigger_ShiftData      <= PortWr[2];
          //Trigger_AudioDeviceP2  <= PortWr[7];
          Trigger_WatchDogReset  <= PortWr[4];
             //<= PortWr[5]; // tone_generator_low_w
             //<= PortWr[6]; // tone_generator_hi_w

	end
        mod_guidedmissle:
        begin 
          // IN0
          GDB0 <= sw[0] | {~m_fire2a,~m_start1,1'b1,1'b1,~m_right2,~m_left2,1'b1,1'b1};
          GDB1 <= sw[1] | {~m_fire1a,~m_start2,1'b1,1'b1,~m_right1,~m_left1,~m_coin1,1'b1};
          // IN2
          GDB2 <= sw[2];
          Trigger_ShiftCount     <= PortWr[1]; // IS THIS WEIRD?
          Trigger_AudioDeviceP1  <= PortWr[3];
          Trigger_ShiftData      <= PortWr[2];
          Trigger_WatchDogReset  <= PortWr[4];
          //<= PortWr[5]; // tone_generator_low_w
          //<= PortWr[6]; // tone_generator_hi_w
	  GDB3 <= ShiftReverse ? SR: S;
        end
        mod_claybust:
        begin 
		    gun_game <= 1;
          // IN0
          GDB1 <= sw[1] | { 1'b0,1'b0,1'b0,1'b0, ~m_start1, ~m_coin1, |claybust_gun_on, |claybust_gun_on};
          GDB2 <=  claybust_gun_pos_lo;
          GDB6 <=  claybust_gun_pos_hi;
          Trigger_ShiftCount     <= PortWr[1];
          Trigger_AudioDeviceP1  <= PortWr[3];
          Trigger_ShiftData      <= PortWr[2];
          Trigger_WatchDogReset  <= PortWr[4];
        end
        mod_gunfight:
	begin
	  WDEnabled <= 1'b0;
          // IN0
          GDB0 <= sw[0] | { m_fire1a,~gunfight_y, m_right1,m_left1,m_down1,m_up1};
          GDB1 <= sw[1] | { m_fire2a,~gunfight_y_2,m_right2,m_left2,m_down2,m_up2};
          GDB2 <= sw[2] | { m_start1,m_coin1, 6'b0};
          Trigger_ShiftCount     <= PortWr[2];
          Trigger_AudioDeviceP1  <= PortWr[1];
          Trigger_ShiftData      <= PortWr[4];
          //Trigger_WatchDogReset  <= PortWr[4];
	end
        mod_indianbattle:
        begin
          landscape<=0;
	  ccw <= 1;
          color_rom_enabled<=1;
          GDB0 <= sw[0];
          GDB1 <= sw[1] | { 1'b1,m_right1,m_left1,m_fire1a, 1'b0,  m_start1,m_start2,~m_coin1};
          GDB2 <= sw[2];
          Trigger_ShiftCount     <= PortWr[2];
          Trigger_AudioDeviceP1  <= PortWr[3];
          Trigger_ShiftData      <= PortWr[4];
          Trigger_AudioDeviceP2  <= PortWr[5];
          Trigger_WatchDogReset  <= PortWr[6];
        end
        mod_lupin:
        begin
          landscape<=0;
	  ccw <= 1;
          GDB0 <= sw[0] | { m_up2,m_left2,m_down2,m_right2,m_fire2a,1'b0,1'b1,1'b1};
          GDB1 <= sw[1] | { m_up1,m_left1,m_down1,m_right1,m_fire1a,m_start1,m_start2,m_coin1};
          GDB2 <= sw[2];
          Trigger_ShiftCount     <= PortWr[2];
          Trigger_AudioDeviceP1  <= PortWr[3];
          Trigger_ShiftData      <= PortWr[4];
          Trigger_AudioDeviceP2  <= PortWr[5];
          Trigger_WatchDogReset  <= PortWr[6];
        end
        mod_m4:
        begin 
          landscape<=1;
	  WDEnabled <= 1'b0;
          // IN0
          GDB0 <= sw[0] | { 1'b1, 1'b1,~m_fire2b,~m_fire2a,~m_down2,1'b1,~m_up2,1'b1};
          GDB1 <= sw[1] | { 1'b1,~m_start2,~m_fire1b,~m_fire1a,~m_down1,~m_start1,~m_up1,~m_coin1};
          GDB2 <= sw[2];
          Trigger_ShiftCount     <= PortWr[1]; // IS THIS WEIRD?
          Trigger_AudioDeviceP1  <= PortWr[3];
          Trigger_ShiftData      <= PortWr[2];
          Trigger_WatchDogReset  <= PortWr[4];
          Trigger_AudioDeviceP2  <= PortWr[5];
	  GDB3 <= ShiftReverse ? SR: S;

        end
        mod_phantom:
        begin
          landscape<=1;
	  GDB0 <= SR;
          GDB1 <= sw[1] | { 1'b1,1'b1,~m_coin1,~m_fire1a,~m_right1,~m_left1,~m_down1,~m_up1};
          GDB2 <= sw[2];
          Trigger_ShiftCount     <= PortWr[1];
          Trigger_ShiftData      <= PortWr[2];
          Trigger_WatchDogReset  <= PortWr[4];
          Trigger_AudioDeviceP1  <= PortWr[5];
          Trigger_AudioDeviceP2  <= PortWr[6];
        end
        mod_polaris:
	begin
          landscape<=0;
	  ccw<=1;
          GDB0 <= sw[0] | { m_up2,m_left2,m_down2,m_right2,m_fire2a,1'b0,1'b0,1'b0};
          GDB1 <= sw[1] | { m_up1,m_left1,m_down1,m_right1,m_fire1a,m_start1,m_start2,m_coin1};
          GDB2 <= sw[2];

          Trigger_ShiftCount     <= PortWr[1];
          Trigger_ShiftData      <= PortWr[3];
          Trigger_WatchDogReset  <= PortWr[5];
          Trigger_AudioDeviceP1  <= PortWr[2];
          Trigger_AudioDeviceP2  <= PortWr[4];
          //<= PortWr[6];

	end
        mod_desertgun:
	begin
          gun_game <= 1;
          landscape <= 1;
          GDB0 <= SR;
          GDB1 <= desert_gun_select ? desert_gun_x[7:0] : desert_gun_y[7:0];
          GDB2 <= sw[2] | { ~m_fire1a,m_coin1, 2'b0, 2'b0, 2'b0};

          Trigger_ShiftCount     <= PortWr[1];
          Trigger_ShiftData      <= PortWr[2];
          Trigger_WatchDogReset  <= PortWr[4];
          Trigger_AudioDeviceP1  <= PortWr[3];
          //<= PortWr[5]; // tone_generator_low_w
          //<= PortWr[6]; // tone_generator_hi_w
          Trigger_AudioDeviceP2  <= PortWr[7];
	end
	mod_seawolf:
	begin
	       gun_game <= 1;
          landscape<=1;
	  WDEnabled <= 1'b0;
          ccw<=0;
          GDB0 <= SR;
	  // IN0
          GDB1 <= sw[0] | { 2'b0, m_fire_a, seawolf_position};
          GDB2 <= sw[1] | { 3'b0,1'b0 /*erase?*/, 2'b0,m_start1,m_coin1};
          Trigger_ShiftData      <= PortWr[3];
          Trigger_ShiftCount     <= PortWr[4];
          //<= PortWr[5];
          //<= PortWr[6];
          //<= PortWr[4];
       end
        mod_yosakdon:
	begin
	  WDEnabled <= 1'b0;
          landscape<=1;
          //GDB0 <= SR;
	  // IN0
          GDB1 <= sw[0] | ~{ 1'b0, m_right,m_left,m_fire_a,1'b0,m_start1, m_start2, m_coin1 };
	  // IN1
          GDB2 <= sw[1] | ~{ 1'b0, m_right,m_left,m_fire_a,1'b0,1'b0,1'b0,1'b0};
	  Trigger_AudioDeviceP1  <= PortWr[3];
          Trigger_AudioDeviceP2  <= PortWr[5];
       end
       mod_spacechaser:
       begin
            landscape<=0;
            ccw<=1;
            color_rom_enabled<=1;
            GDB0 <= sw[0] | { 1'b0, 1'b0,1'b0,  m_fire2a,  m_right2,m_down2,m_left2,m_up2};
            GDB1 <= sw[1] | { m_coin1,m_start1,m_start2,m_fire_a,m_right,m_down,m_left,m_up};
            GDB2 <= sw[2];
       end
       mod_steelworker:
       begin
	  WDEnabled <= 1'b0;
           GDB0 <= 0;
	   GDB1 <= sw[1] |{ ~m_fire1b, m_right,m_left,m_fire1a,1'b0,m_start1,m_start2, ~m_coin1};
	   GDB2 <= sw[2] |{ ~m_fire2b, m_right2, m_left2 , m_fire2a,1'b0,1'b0, 1'b0,1'b0} ;
           Trigger_ShiftCount     <= PortWr[2];
          //Trigger_AudioDeviceP1  <= PortWr[2];
          Trigger_ShiftData      <= PortWr[4];
          //Trigger_AudioDeviceP2  <= PortWr[5];
          //Trigger_WatchDogReset  <= PortWr[7];
       end
      endcase
end

wire [15:0] color_prom_addr;
wire [7:0]  color_prom_out;
wire [15:0]RAB;
wire [15:0]AD;
wire [7:0]RDB;
wire [7:0]RWD;
wire [7:0]IB;
wire [5:0]SoundCtrl3;
wire [5:0]SoundCtrl5;
wire Rst_n_s;
wire RWE_n;
wire Video;
wire HSync;
wire VSync;
wire CPU_RW_n;

invaderst invaderst(
        .Rst_n(~(reset)),
        .Clk(clk_sys),
        .ENA(),
		  
        .GDB0(GDB0),
        .GDB1(GDB1),
        .GDB2(GDB2),
        .GDB3(GDB3),
        .GDB4(GDB4),
        .GDB5(GDB5),
        .GDB6(GDB6),

	.WD_Enabled(WDEnabled),

        .RDB(RDB),
        .IB(IB),
        .RWD(RWD),
        .RAB(RAB),
        .AD(AD),
        .SoundCtrl3(SoundCtrl3),
        .SoundCtrl5(SoundCtrl5),
        .Rst_n_s(Rst_n_s),
        .RWE_n(RWE_n),
        .Video(Video),
		  .CPU_RW_n(CPU_RW_n),

	.color_prom_addr(color_prom_addr),
	.color_prom_out(color_prom_out),
        .O_VIDEO_R(r),
        .O_VIDEO_G(g),
        .O_VIDEO_B(b),
        //.HBLANK(hblank),
        //.VBLANK(vblank),
        .Overlay(~status[8]),
	.OverlayTest(status[9]),

        .HSync(HSync),
        .VSync(VSync),


        .Trigger_ShiftCount(Trigger_ShiftCount),
        .Trigger_ShiftData(Trigger_ShiftData),
        .Trigger_AudioDeviceP1(Trigger_AudioDeviceP1),
        .Trigger_AudioDeviceP2(Trigger_AudioDeviceP2),
        .Trigger_WatchDogReset(Trigger_WatchDogReset),

        .PortWr(PortWr),
        .S(S),
        .ShiftReverse(ShiftReverse),

	.mod_vortex(mod==mod_vortex)
        );
invaders_memory invaders_memory (
        .Clock(clk_sys),
        .RW_n(RWE_n),
		  .CPU_RW_n(CPU_RW_n),
        .Addr(AD),
        .Ram_Addr(RAB),
        .Ram_out(RDB),
        .Ram_in(RWD),
        .Rom_out(IB),
	.color_prom_out(color_prom_out),
	.color_prom_addr(color_prom_addr),

	.dn_addr(ioctl_addr[15:0]),
	.dn_data(ioctl_dout),
	.dn_wr(ioctl_wr&ioctl_index==0),
	.mod_vortex(mod==mod_vortex),
	.mod_attackforce(mod==mod_attackforce),
	.mod_cosmo(mod==mod_cosmo)
        );

invaders_audio invaders_audio (
        .Clk(clk_sys),
        .S1(SoundCtrl3),
        .S2(SoundCtrl5),
        .Aud(inv_audio_data)
        );

zap_audio zap_audio (
        .Clk(clk_sys),
        .S1(SoundCtrl3),
        .S2(SoundCtrl5),
        .Aud(zap_audio_data)
        );

invaders_blank invaders_blank (
        .CLK(clk_sys),
        .Rst_n_s(Rst_n_s),
        .HSync(HSync),
        .VSync(VSync),
        .O_HBLANK(hblank),
        .O_VBLANK(vblank)
	);




wire bg_download = ioctl_download && (ioctl_index == 2);

reg [7:0] ioctl_dout_r;
always @(posedge clk_sys) if(ioctl_wr & ~ioctl_addr[0]) ioctl_dout_r <= ioctl_dout;

wire [31:0] pic_data;
sdram sdram
(
	.*,

	.init(~pll_locked),
	.clk(clk_mem),
	.ch1_addr(bg_download ? ioctl_addr[24:1] : pic_addr),
	.ch1_dout(pic_data),
	.ch1_din({ioctl_dout, ioctl_dout_r}),
	.ch1_req(bg_download ? (ioctl_wr & ioctl_addr[0]) : pic_req),
	.ch1_rnw(~bg_download)
);

reg        pic_req;
reg [24:1] pic_addr;
reg  [7:0] bg_r,bg_g,bg_b,bg_a;
always @(posedge clk_40) begin
	reg old_vs;
	reg use_bg = 0;
	
	if(bg_download && sdram_sz[2:0]) use_bg <= 1;

	pic_req <= 0;

	if(use_bg) begin
		if(ce_pix) begin
			old_vs <= VSync;
			{bg_a,bg_b,bg_g,bg_r} <= pic_data;
			if(~(hblank|vblank)) begin
				pic_addr <= pic_addr + 2'd2;
				pic_req <= 1;
			end
			
			if(~old_vs & VSync) begin
				pic_addr <= 0;
				pic_req <= 1;
			end
		end
	end
	else begin
		{bg_a,bg_b,bg_g,bg_r} <= 0;
	end
end

wire [1:0] gun_mode = status[12:11];
wire [1:0] gun_cross_size = status[14:13];
wire       gun_target;
wire [7:0] gun_x, gun_y;
reg        gun_game = 0;

virtualgun virtualgun
(
	.CLK(clk_40),
	
	.MOUSE(ps2_mouse),
	.MOUSE_XY(gun_mode[1]),
	.JOY_X(!gun_mode ? joya[7:0] : joya2[7:0]),
	.JOY_Y(!gun_mode ? joya[15:8] : joya2[15:8]),
	.JOY(!gun_mode ? joy1 : joy2),

	.HDE(~hblank),
	.VDE(~vblank),
	.CE_PIX(ce_pix),

	.SIZE(gun_cross_size),

	.TARGET(gun_target),
	.X_OUT(gun_x),
	.Y_OUT(gun_y)
);

endmodule
