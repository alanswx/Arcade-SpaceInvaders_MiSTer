library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity cv18_35 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of cv18_35 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"CD",X"B4",X"19",X"06",X"20",X"CD",X"F0",X"18",X"CD",X"2D",X"16",X"CD",X"82",X"15",X"CD",
		X"08",X"16",X"CD",X"7A",X"09",X"3A",X"82",X"20",X"A7",X"CA",X"DE",X"09",X"CD",X"21",X"17",X"CD",
		X"21",X"09",X"CD",X"BC",X"08",X"CD",X"4A",X"17",X"CD",X"48",X"0A",X"CA",X"33",X"08",X"06",X"04",
		X"CD",X"F0",X"18",X"CD",X"91",X"17",X"D3",X"06",X"CD",X"14",X"18",X"C3",X"09",X"08",X"11",X"BA",
		X"1A",X"CD",X"DF",X"08",X"06",X"98",X"DB",X"01",X"0F",X"0F",X"DA",X"54",X"08",X"0F",X"DA",X"7F",
		X"07",X"C3",X"66",X"07",X"3E",X"01",X"C3",X"82",X"07",X"CD",X"02",X"02",X"C3",X"FE",X"07",X"3A",
		X"08",X"20",X"47",X"2A",X"09",X"20",X"EB",X"C3",X"6A",X"08",X"3A",X"67",X"20",X"67",X"2E",X"FC",
		X"C9",X"21",X"11",X"2B",X"11",X"70",X"1B",X"0E",X"0E",X"CD",X"DF",X"08",X"3A",X"67",X"20",X"0F",
		X"3E",X"1C",X"21",X"11",X"37",X"D4",X"EB",X"08",X"3E",X"B0",X"32",X"C0",X"20",X"3A",X"C0",X"20",
		X"A7",X"C8",X"E6",X"04",X"C2",X"A0",X"08",X"CD",X"B9",X"09",X"CD",X"18",X"19",X"C3",X"8D",X"08",
		X"06",X"28",X"21",X"1C",X"27",X"3A",X"67",X"20",X"0F",X"DA",X"AF",X"08",X"21",X"1C",X"39",X"CD",
		X"84",X"14",X"C3",X"8D",X"08",X"DB",X"02",X"E6",X"03",X"C6",X"03",X"C9",X"3A",X"82",X"20",X"FE",
		X"09",X"D0",X"3E",X"FB",X"32",X"7E",X"20",X"C9",X"3E",X"02",X"32",X"FB",X"21",X"32",X"FB",X"22",
		X"3A",X"CE",X"20",X"A7",X"C0",X"21",X"1C",X"39",X"06",X"28",X"C3",X"84",X"14",X"0E",X"03",X"1A",
		X"D5",X"CD",X"EB",X"08",X"D1",X"13",X"0D",X"C2",X"DF",X"08",X"C9",X"11",X"00",X"1E",X"E5",X"26",
		X"00",X"6F",X"29",X"29",X"29",X"19",X"EB",X"E1",X"06",X"08",X"D3",X"06",X"C3",X"15",X"14",X"3A",
		X"09",X"20",X"FE",X"78",X"D0",X"2A",X"91",X"20",X"7D",X"B4",X"C2",X"15",X"09",X"21",X"00",X"06",
		X"3E",X"01",X"32",X"83",X"20",X"2B",X"22",X"91",X"20",X"C9",X"CD",X"26",X"16",X"2E",X"FF",X"7E",
		X"C9",X"CD",X"FA",X"18",X"2B",X"2B",X"7E",X"A7",X"C8",X"06",X"15",X"DB",X"02",X"E6",X"08",X"CA",
		X"34",X"09",X"06",X"10",X"CD",X"3D",X"17",X"B8",X"D8",X"CD",X"1A",X"09",X"34",X"7E",X"F5",X"21",
		X"01",X"25",X"24",X"24",X"3D",X"C2",X"42",X"09",X"06",X"10",X"11",X"60",X"1C",X"CD",X"15",X"14",
		X"F1",X"3C",X"CD",X"71",X"1A",X"CD",X"FA",X"18",X"2B",X"2B",X"36",X"00",X"3E",X"FF",X"32",X"99",
		X"20",X"06",X"10",X"C3",X"F0",X"18",X"21",X"A0",X"1D",X"FE",X"02",X"D8",X"23",X"FE",X"04",X"D8",
		X"23",X"C9",X"CD",X"9C",X"09",X"3E",X"1A",X"C3",X"EB",X"08",X"CD",X"B9",X"09",X"3A",X"F1",X"20",
		X"A7",X"C8",X"AF",X"32",X"F1",X"20",X"E5",X"2A",X"F2",X"20",X"EB",X"E1",X"7E",X"83",X"27",X"77",
		X"5F",X"23",X"7E",X"8A",X"27",X"77",X"57",X"23",X"7E",X"23",X"66",X"6F",X"7A",X"CD",X"A1",X"09",
		X"7B",X"D5",X"F5",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"CD",X"B4",X"09",X"F1",X"E6",X"0F",X"CD",
		X"B4",X"09",X"D1",X"C9",X"C6",X"1A",X"C3",X"EB",X"08",X"3A",X"67",X"20",X"0F",X"21",X"F8",X"20",
		X"D8",X"21",X"FC",X"20",X"C9",X"21",X"02",X"24",X"36",X"00",X"23",X"7D",X"E6",X"1F",X"FE",X"1C",
		X"DA",X"D7",X"09",X"11",X"06",X"00",X"19",X"7C",X"FE",X"40",X"DA",X"C8",X"09",X"C9",X"CD",X"28",
		X"0A",X"AF",X"32",X"E9",X"20",X"CD",X"C5",X"09",X"3A",X"67",X"20",X"F5",X"CD",X"CC",X"01",X"F1",
		X"32",X"67",X"20",X"67",X"E5",X"2E",X"FE",X"7E",X"E6",X"07",X"3C",X"77",X"21",X"A2",X"1D",X"23",
		X"3D",X"C2",X"FF",X"09",X"7E",X"E1",X"2E",X"FC",X"77",X"23",X"36",X"38",X"7C",X"0F",X"DA",X"1F",
		X"0A",X"3E",X"21",X"32",X"98",X"20",X"CD",X"DD",X"01",X"CD",X"A2",X"01",X"C3",X"EE",X"07",X"CD",
		X"D7",X"01",X"CD",X"A8",X"01",X"C3",X"EE",X"07",X"CD",X"48",X"0A",X"C2",X"41",X"0A",X"3E",X"30",
		X"32",X"C0",X"20",X"3A",X"C0",X"20",X"A7",X"C8",X"CD",X"48",X"0A",X"CA",X"33",X"0A",X"CD",X"5B",
		X"14",X"CD",X"48",X"0A",X"C2",X"41",X"0A",X"C9",X"3A",X"15",X"20",X"FE",X"FF",X"C9",X"3A",X"EF",
		X"20",X"A7",X"CA",X"6B",X"0A",X"48",X"06",X"08",X"CD",X"F0",X"18",X"41",X"78",X"CD",X"66",X"09",
		X"7E",X"21",X"F3",X"20",X"36",X"00",X"2B",X"77",X"2B",X"36",X"01",X"21",X"62",X"20",X"C9",X"3E",
		X"02",X"32",X"C1",X"20",X"D3",X"06",X"3A",X"CB",X"20",X"A7",X"CA",X"74",X"0A",X"AF",X"32",X"C1",
		X"20",X"C9",X"D5",X"1A",X"CD",X"EB",X"08",X"D1",X"3E",X"07",X"32",X"C0",X"20",X"3A",X"C0",X"20",
		X"3D",X"C2",X"8D",X"0A",X"13",X"0D",X"C2",X"82",X"0A",X"C9",X"21",X"50",X"20",X"C3",X"33",X"02",
		X"3E",X"40",X"C3",X"C6",X"0A",X"3E",X"80",X"C3",X"C6",X"0A",X"E1",X"C3",X"72",X"00",X"3A",X"C1",
		X"20",X"0F",X"DA",X"AA",X"0A",X"0F",X"DA",X"75",X"18",X"0F",X"DA",X"9A",X"0A",X"C9",X"21",X"14",
		X"2B",X"0E",X"0F",X"C3",X"82",X"0A",X"32",X"C0",X"20",X"3A",X"C0",X"20",X"A7",X"C2",X"C9",X"0A",
		X"C9",X"21",X"C2",X"20",X"06",X"0C",X"C3",X"14",X"1A",X"31",X"00",X"24",X"06",X"00",X"CD",X"CE",
		X"01",X"CD",X"3D",X"19",X"3E",X"08",X"32",X"CF",X"20",X"AF",X"D3",X"03",X"D3",X"05",X"CD",X"69",
		X"19",X"FB",X"CD",X"A0",X"0A",X"3A",X"EC",X"20",X"A7",X"21",X"17",X"30",X"0E",X"04",X"C2",X"E7",
		X"0B",X"11",X"FA",X"1C",X"CD",X"82",X"0A",X"11",X"AF",X"1D",X"CD",X"BE",X"0A",X"CD",X"A0",X"0A",
		X"CD",X"25",X"18",X"CD",X"A5",X"0A",X"3A",X"EC",X"20",X"A7",X"C2",X"49",X"0B",X"11",X"95",X"1A",
		X"CD",X"D1",X"0A",X"CD",X"6F",X"0A",X"11",X"B0",X"1B",X"CD",X"D1",X"0A",X"CD",X"6F",X"0A",X"CD",
		X"A0",X"0A",X"11",X"C9",X"1F",X"CD",X"D1",X"0A",X"CD",X"6F",X"0A",X"CD",X"A0",X"0A",X"21",X"F7",
		X"33",X"06",X"0A",X"CD",X"84",X"14",X"CD",X"A5",X"0A",X"CD",X"C5",X"09",X"3A",X"FF",X"21",X"A7",
		X"C2",X"5C",X"0B",X"CD",X"B5",X"08",X"32",X"FF",X"21",X"CD",X"65",X"1A",X"CD",X"CC",X"01",X"CD",
		X"A8",X"01",X"CD",X"D7",X"01",X"CD",X"02",X"02",X"3E",X"01",X"32",X"C1",X"20",X"CD",X"B7",X"01",
		X"CD",X"2D",X"16",X"CD",X"F0",X"0B",X"D3",X"06",X"CD",X"48",X"0A",X"CA",X"70",X"0B",X"AF",X"32",
		X"25",X"20",X"CD",X"48",X"0A",X"C2",X"82",X"0B",X"AF",X"32",X"C1",X"20",X"CD",X"A0",X"0A",X"CD",
		X"6F",X"19",X"0E",X"0C",X"21",X"11",X"2C",X"11",X"90",X"1F",X"CD",X"DF",X"08",X"3A",X"EC",X"20",
		X"FE",X"00",X"C2",X"AD",X"0B",X"21",X"11",X"33",X"3E",X"02",X"CD",X"EB",X"08",X"01",X"9C",X"1F",
		X"CD",X"63",X"18",X"CD",X"59",X"18",X"DB",X"02",X"07",X"DA",X"C2",X"0B",X"01",X"A0",X"1F",X"CD",
		X"47",X"18",X"CD",X"A5",X"0A",X"3A",X"EC",X"20",X"FE",X"00",X"C2",X"D9",X"0B",X"11",X"D5",X"1F",
		X"CD",X"D1",X"0A",X"CD",X"6F",X"0A",X"CD",X"A8",X"18",X"21",X"EC",X"20",X"7E",X"3C",X"E6",X"01",
		X"77",X"CD",X"C5",X"09",X"C3",X"E4",X"0A",X"11",X"AB",X"1D",X"CD",X"82",X"0A",X"C3",X"0A",X"0B",
		X"CD",X"82",X"15",X"C3",X"7D",X"19",X"13",X"00",X"08",X"13",X"0E",X"26",X"02",X"0E",X"0F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
